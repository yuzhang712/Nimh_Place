# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405300513        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Tue, 3 Jun 2014, 13:07:07.
# Main process id is 12480.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2_X1_8T
  CLASS core ;
  FOREIGN AND2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.4639 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0847 0.078 0.35 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.076 0.334 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.108 0.1419 0.1267 ;
        RECT 0.114 0.1267 0.1419 0.2853 ;
        RECT 0.114 0.2853 0.1419 0.3627 ;
        RECT 0.1419 0.108 0.242 0.1267 ;
        RECT 0.242 0.108 0.27 0.1267 ;
        RECT 0.242 0.1267 0.27 0.2853 ;
      LAYER M1 ;
        RECT 0.114 0.108 0.1419 0.1267 ;
        RECT 0.114 0.1267 0.1419 0.2853 ;
        RECT 0.114 0.2853 0.1419 0.3627 ;
        RECT 0.1419 0.108 0.242 0.1267 ;
        RECT 0.242 0.108 0.27 0.1267 ;
        RECT 0.242 0.1267 0.27 0.2853 ;
  END
END AND2_X1_8T

MACRO AND2_X2_8T
  CLASS core ;
  FOREIGN AND2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1653 0.083 0.3467 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.0427 0.306 0.0867 ;
        RECT 0.302 0.4253 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.0867 ;
        RECT 0.306 0.0867 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.3827 0.082 0.4013 ;
        RECT 0.082 0.1107 0.242 0.1293 ;
        RECT 0.082 0.3827 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.1293 ;
        RECT 0.242 0.1293 0.27 0.3827 ;
        RECT 0.242 0.3827 0.27 0.4013 ;
      LAYER M1 ;
        RECT 0.054 0.3827 0.082 0.4013 ;
        RECT 0.082 0.1107 0.242 0.1293 ;
        RECT 0.082 0.3827 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.1293 ;
        RECT 0.242 0.1293 0.27 0.3827 ;
        RECT 0.242 0.3827 0.27 0.4013 ;
  END
END AND2_X2_8T

MACRO AND3_X1_8T
  CLASS core ;
  FOREIGN AND3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1729 0.128 0.211 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.128 0.08 0.384 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.076 0.462 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.079 0.0667 0.238 0.066732 ;
        RECT 0.054 0.4207 0.274 0.4393 ;
        RECT 0.274 0.0633 0.37 0.0913 ;
        RECT 0.274 0.4207 0.37 0.4393 ;
        RECT 0.37 0.0633 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4393 ;
      LAYER M1 ;
        RECT 0.079 0.0667 0.238 0.066732 ;
        RECT 0.054 0.4207 0.274 0.4393 ;
        RECT 0.274 0.0633 0.37 0.0913 ;
        RECT 0.274 0.4207 0.37 0.4393 ;
        RECT 0.37 0.0633 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4393 ;
  END
END AND3_X1_8T

MACRO AND3_X2_8T
  CLASS core ;
  FOREIGN AND3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.2133 0.206 0.342 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1707 0.083 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2013 0.27 0.358 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.0427 0.37 0.1047 ;
        RECT 0.366 0.4253 0.37 0.4693 ;
        RECT 0.37 0.0427 0.398 0.1047 ;
        RECT 0.37 0.1047 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.048 0.08 0.104 ;
        RECT 0.048 0.104 0.08 0.1253 ;
        RECT 0.08 0.104 0.298 0.1253 ;
        RECT 0.054 0.3873 0.146 0.4087 ;
        RECT 0.146 0.1493 0.306 0.168 ;
        RECT 0.146 0.3873 0.306 0.4087 ;
        RECT 0.306 0.1493 0.334 0.168 ;
        RECT 0.306 0.168 0.334 0.3873 ;
        RECT 0.306 0.3873 0.334 0.4087 ;
      LAYER M1 ;
        RECT 0.048 0.048 0.08 0.104 ;
        RECT 0.048 0.104 0.08 0.1253 ;
        RECT 0.08 0.104 0.298 0.1253 ;
        RECT 0.054 0.3873 0.146 0.4087 ;
        RECT 0.146 0.1493 0.306 0.168 ;
        RECT 0.146 0.3873 0.306 0.4087 ;
        RECT 0.306 0.1493 0.334 0.168 ;
        RECT 0.306 0.168 0.334 0.3873 ;
        RECT 0.306 0.3873 0.334 0.4087 ;
  END
END AND3_X2_8T

MACRO AND4_X1_8T
  CLASS core ;
  FOREIGN AND4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.128 0.272 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.3413 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.076 0.526 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.424 0.338 0.4453 ;
        RECT 0.338 0.0667 0.434 0.066732 ;
        RECT 0.338 0.424 0.434 0.4453 ;
        RECT 0.434 0.0667 0.462 0.066732 ;
        RECT 0.434 0.088 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
        RECT 0.1409 0.066 0.298 0.098 ;
      LAYER M1 ;
        RECT 0.082 0.424 0.338 0.4453 ;
        RECT 0.338 0.0667 0.434 0.066732 ;
        RECT 0.338 0.424 0.434 0.4453 ;
        RECT 0.434 0.0667 0.462 0.066732 ;
        RECT 0.434 0.088 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
        RECT 0.1409 0.066 0.298 0.098 ;
  END
END AND4_X1_8T

MACRO AND4_X2_8T
  CLASS core ;
  FOREIGN AND4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1607 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.128 0.27 0.3847 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.3847 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.3847 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.064 0.526 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0667419 0.0667 0.298 0.066732 ;
        RECT 0.082 0.424 0.342 0.4453 ;
        RECT 0.342 0.11 0.434 0.1313 ;
        RECT 0.342 0.424 0.434 0.4453 ;
        RECT 0.434 0.11 0.462 0.1313 ;
        RECT 0.434 0.1313 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
      LAYER M1 ;
        RECT 0.0667419 0.0667 0.298 0.066732 ;
        RECT 0.082 0.424 0.342 0.4453 ;
        RECT 0.342 0.11 0.434 0.1313 ;
        RECT 0.342 0.424 0.434 0.4453 ;
        RECT 0.434 0.11 0.462 0.1313 ;
        RECT 0.434 0.1313 0.462 0.424 ;
        RECT 0.434 0.424 0.462 0.4453 ;
  END
END AND4_X2_8T

MACRO ANTENNA_8T
  CLASS core ;
  FOREIGN ANTENNA_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
END ANTENNA_8T

MACRO AOI21_X1_8T
  CLASS core ;
  FOREIGN AOI21_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.128 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0893 0.078 0.3413 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.3413 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.066714 0.0667 0.0667419 0.066732 ;
        RECT 0.114 0.088 0.1419 0.3573 ;
        RECT 0.0667419 0.0667 0.306 0.066732 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3867 0.08 0.408 ;
        RECT 0.048 0.408 0.08 0.4693 ;
        RECT 0.08 0.3867 0.298 0.408 ;
      LAYER M1 ;
        RECT 0.048 0.3867 0.08 0.408 ;
        RECT 0.048 0.408 0.08 0.4693 ;
        RECT 0.08 0.3867 0.298 0.408 ;
  END
END AOI21_X1_8T

MACRO AOI21_X2_8T
  CLASS core ;
  FOREIGN AOI21_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.2013 0.398 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1533 0.27 0.172 ;
        RECT 0.242 0.172 0.27 0.2987 ;
        RECT 0.242 0.2987 0.27 0.3413 ;
        RECT 0.27 0.1533 0.493 0.172 ;
        RECT 0.493 0.1533 0.531 0.172 ;
        RECT 0.493 0.172 0.531 0.2987 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.2987 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.077 0.1107 0.178 0.1293 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.326 ;
        RECT 0.178 0.326 0.206 0.3806 ;
        RECT 0.178 0.3806 0.206 0.3993 ;
        RECT 0.206 0.1107 0.43 0.1293 ;
        RECT 0.206 0.3806 0.43 0.3993 ;
        RECT 0.43 0.3806 0.434 0.3993 ;
        RECT 0.434 0.326 0.462 0.3806 ;
        RECT 0.434 0.3806 0.462 0.3993 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3667 0.08 0.4233 ;
        RECT 0.048 0.4233 0.08 0.446 ;
        RECT 0.08 0.4233 0.498 0.446 ;
        RECT 0.498 0.344 0.526 0.3667 ;
        RECT 0.498 0.3667 0.526 0.4233 ;
        RECT 0.498 0.4233 0.526 0.446 ;
        RECT 0.146 0.0679 0.535 0.0867 ;
      LAYER M1 ;
        RECT 0.048 0.3667 0.08 0.4233 ;
        RECT 0.048 0.4233 0.08 0.446 ;
        RECT 0.08 0.4233 0.498 0.446 ;
        RECT 0.498 0.344 0.526 0.3667 ;
        RECT 0.498 0.3667 0.526 0.4233 ;
        RECT 0.498 0.4233 0.526 0.446 ;
        RECT 0.146 0.0679 0.535 0.0867 ;
  END
END AOI21_X2_8T

MACRO AOI22_X1_8T
  CLASS core ;
  FOREIGN AOI22_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.128 0.27 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.3233 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.132 0.1419 0.384 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.0679 0.306 0.0867 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.0867 0.334 0.388 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.42 0.37 0.4493 ;
        RECT 0.37 0.3687 0.398 0.42 ;
        RECT 0.37 0.42 0.398 0.4493 ;
      LAYER M1 ;
        RECT 0.082 0.42 0.37 0.4493 ;
        RECT 0.37 0.3687 0.398 0.42 ;
        RECT 0.37 0.42 0.398 0.4493 ;
  END
END AOI22_X1_8T

MACRO AOI22_X2_8T
  CLASS core ;
  FOREIGN AOI22_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.1827 0.462 0.2013 ;
        RECT 0.434 0.2013 0.462 0.326 ;
        RECT 0.434 0.326 0.462 0.3413 ;
        RECT 0.462 0.1827 0.654 0.2013 ;
        RECT 0.654 0.1827 0.6899 0.2013 ;
        RECT 0.6899 0.1827 0.718 0.2013 ;
        RECT 0.6899 0.2013 0.718 0.326 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.2467 0.59 0.3413 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.204 0.204 0.334 0.3507 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1613 0.078 0.3413 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.133342 0.1333 0.13337 0.133328 ;
        RECT 0.242 0.152 0.27 0.1527 ;
        RECT 0.242 0.1527 0.27 0.2133 ;
        RECT 0.13337 0.1333 0.362 0.133328 ;
        RECT 0.362 0.1333 0.37 0.133328 ;
        RECT 0.37 0.1333 0.398 0.133328 ;
        RECT 0.37 0.152 0.398 0.1527 ;
        RECT 0.37 0.1527 0.398 0.2133 ;
        RECT 0.37 0.2133 0.398 0.3087 ;
        RECT 0.37 0.3087 0.398 0.3786 ;
        RECT 0.37 0.3786 0.398 0.4013 ;
        RECT 0.398 0.1333 0.626 0.133328 ;
        RECT 0.398 0.152 0.626 0.1527 ;
        RECT 0.398 0.3786 0.626 0.4013 ;
        RECT 0.626 0.1333 0.654 0.133328 ;
        RECT 0.626 0.152 0.654 0.1527 ;
        RECT 0.626 0.3087 0.654 0.3786 ;
        RECT 0.626 0.3786 0.654 0.4013 ;
        RECT 0.654 0.1333 0.6899 0.133328 ;
        RECT 0.654 0.152 0.6899 0.1527 ;
        RECT 0.6899 0.064 0.718 0.1333 ;
        RECT 0.6899 0.1333 0.718 0.133328 ;
        RECT 0.6899 0.152 0.718 0.1527 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.406 0.088 0.626 0.1093 ;
        RECT 0.626 0.048 0.654 0.088 ;
        RECT 0.626 0.088 0.654 0.1093 ;
        RECT 0.077 0.4253 0.6899 0.444 ;
        RECT 0.6899 0.3713 0.718 0.4253 ;
        RECT 0.6899 0.4253 0.718 0.444 ;
        RECT 0.0859 0.0579 0.362 0.0967 ;
      LAYER M1 ;
        RECT 0.406 0.088 0.626 0.1093 ;
        RECT 0.626 0.048 0.654 0.088 ;
        RECT 0.626 0.088 0.654 0.1093 ;
        RECT 0.077 0.4253 0.6899 0.444 ;
        RECT 0.6899 0.3713 0.718 0.4253 ;
        RECT 0.6899 0.4253 0.718 0.444 ;
        RECT 0.0859 0.0579 0.362 0.0967 ;
  END
END AOI22_X2_8T

MACRO BUF_X1_8T
  CLASS core ;
  FOREIGN BUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.076 0.272 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1429 0.5307 ;
        RECT 0.1429 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.2853 0.115 0.304 ;
        RECT 0.114 0.304 0.115 0.372 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.2853 ;
        RECT 0.115 0.2853 0.1419 0.304 ;
        RECT 0.115 0.304 0.1419 0.372 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.2853 ;
        RECT 0.1419 0.2853 0.1429 0.304 ;
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.2853 0.115 0.304 ;
        RECT 0.114 0.304 0.115 0.372 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.2853 ;
        RECT 0.115 0.2853 0.1419 0.304 ;
        RECT 0.115 0.304 0.1419 0.372 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.2853 ;
        RECT 0.1419 0.2853 0.1429 0.304 ;
  END
END BUF_X1_8T

MACRO BUF_X2_8T
  CLASS core ;
  FOREIGN BUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.178 0.078 0.3413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.402 0.177 0.4693 ;
        RECT 0.177 0.048 0.178 0.088 ;
        RECT 0.177 0.402 0.178 0.4693 ;
        RECT 0.178 0.048 0.206 0.088 ;
        RECT 0.178 0.088 0.206 0.402 ;
        RECT 0.178 0.402 0.206 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.042 0.3707 0.05 0.3893 ;
        RECT 0.042 0.3893 0.05 0.4573 ;
        RECT 0.05 0.064 0.078 0.128 ;
        RECT 0.05 0.128 0.078 0.1467 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4573 ;
        RECT 0.078 0.128 0.0859 0.1467 ;
        RECT 0.078 0.3707 0.0859 0.3893 ;
        RECT 0.078 0.3893 0.0859 0.4573 ;
        RECT 0.0859 0.128 0.114 0.1467 ;
        RECT 0.0859 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
      LAYER M1 ;
        RECT 0.042 0.3707 0.05 0.3893 ;
        RECT 0.042 0.3893 0.05 0.4573 ;
        RECT 0.05 0.064 0.078 0.128 ;
        RECT 0.05 0.128 0.078 0.1467 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4573 ;
        RECT 0.078 0.128 0.0859 0.1467 ;
        RECT 0.078 0.3707 0.0859 0.3893 ;
        RECT 0.078 0.3893 0.0859 0.4573 ;
        RECT 0.0859 0.128 0.114 0.1467 ;
        RECT 0.0859 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
  END
END BUF_X2_8T

MACRO BUF_X4_8T
  CLASS core ;
  FOREIGN BUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1613 0.206 0.3507 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.0679 0.21 0.0867 ;
        RECT 0.21 0.0679 0.27 0.0867 ;
        RECT 0.21 0.4253 0.27 0.444 ;
        RECT 0.27 0.0679 0.368 0.0867 ;
        RECT 0.27 0.4253 0.368 0.444 ;
        RECT 0.368 0.0679 0.4 0.0867 ;
        RECT 0.368 0.0867 0.4 0.4253 ;
        RECT 0.368 0.4253 0.4 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.027 0.1107 0.0859 0.132 ;
        RECT 0.0859 0.1107 0.242 0.132 ;
        RECT 0.0859 0.3799 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.132 ;
        RECT 0.242 0.132 0.27 0.3799 ;
        RECT 0.242 0.3799 0.27 0.4013 ;
      LAYER M1 ;
        RECT 0.027 0.1107 0.0859 0.132 ;
        RECT 0.0859 0.1107 0.242 0.132 ;
        RECT 0.0859 0.3799 0.242 0.4013 ;
        RECT 0.242 0.1107 0.27 0.132 ;
        RECT 0.242 0.132 0.27 0.3799 ;
        RECT 0.242 0.3799 0.27 0.4013 ;
  END
END BUF_X4_8T

MACRO BUF_X8_8T
  CLASS core ;
  FOREIGN BUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.244 ;
        RECT 0.05 0.244 0.078 0.2653 ;
        RECT 0.05 0.2653 0.078 0.3413 ;
        RECT 0.078 0.244 0.298 0.2653 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.0679 0.7 0.0867 ;
        RECT 0.338 0.4253 0.7 0.444 ;
        RECT 0.7 0.0679 0.754 0.0867 ;
        RECT 0.7 0.4253 0.754 0.444 ;
        RECT 0.754 0.0679 0.782 0.0867 ;
        RECT 0.754 0.0867 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.7 0.5307 ;
        RECT 0.7 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.099 0.0653 0.114 0.124 ;
        RECT 0.099 0.124 0.114 0.1427 ;
        RECT 0.114 0.0653 0.1419 0.124 ;
        RECT 0.114 0.124 0.1419 0.1427 ;
        RECT 0.114 0.3513 0.1419 0.3887 ;
        RECT 0.114 0.3887 0.1419 0.4467 ;
        RECT 0.1419 0.0653 0.157 0.124 ;
        RECT 0.1419 0.124 0.157 0.1427 ;
        RECT 0.1419 0.3513 0.157 0.3887 ;
        RECT 0.157 0.124 0.354 0.1427 ;
        RECT 0.157 0.3513 0.354 0.3887 ;
        RECT 0.354 0.124 0.382 0.1427 ;
        RECT 0.354 0.1427 0.382 0.2273 ;
        RECT 0.354 0.2273 0.382 0.246 ;
        RECT 0.354 0.246 0.382 0.3513 ;
        RECT 0.354 0.3513 0.382 0.3887 ;
        RECT 0.382 0.2273 0.7 0.246 ;
      LAYER M1 ;
        RECT 0.099 0.0653 0.114 0.124 ;
        RECT 0.099 0.124 0.114 0.1427 ;
        RECT 0.114 0.0653 0.1419 0.124 ;
        RECT 0.114 0.124 0.1419 0.1427 ;
        RECT 0.114 0.3513 0.1419 0.3887 ;
        RECT 0.114 0.3887 0.1419 0.4467 ;
        RECT 0.1419 0.0653 0.157 0.124 ;
        RECT 0.1419 0.124 0.157 0.1427 ;
        RECT 0.1419 0.3513 0.157 0.3887 ;
        RECT 0.157 0.124 0.354 0.1427 ;
        RECT 0.157 0.3513 0.354 0.3887 ;
        RECT 0.354 0.124 0.382 0.1427 ;
        RECT 0.354 0.1427 0.382 0.2273 ;
        RECT 0.354 0.2273 0.382 0.246 ;
        RECT 0.354 0.246 0.382 0.3513 ;
        RECT 0.354 0.3513 0.382 0.3887 ;
        RECT 0.382 0.2273 0.7 0.246 ;
  END
END BUF_X8_8T

MACRO BUF_X12_8T
  CLASS core ;
  FOREIGN BUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.1573 0.08 0.244 ;
        RECT 0.048 0.244 0.08 0.2653 ;
        RECT 0.048 0.2653 0.08 0.3433 ;
        RECT 0.08 0.244 0.426 0.2653 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.0679 1.07 0.0867 ;
        RECT 0.466 0.4253 1.07 0.444 ;
        RECT 1.07 0.0679 1.1359 0.0867 ;
        RECT 1.07 0.4253 1.1359 0.444 ;
        RECT 1.1359 0.0679 1.168 0.0867 ;
        RECT 1.1359 0.0867 1.168 0.4253 ;
        RECT 1.1359 0.4253 1.168 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.07 0.5307 ;
        RECT 1.07 0.4933 1.29 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.29 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.098 0.3673 0.112 0.3887 ;
        RECT 0.098 0.3887 0.112 0.4467 ;
        RECT 0.112 0.0653 0.144 0.1233 ;
        RECT 0.112 0.1233 0.144 0.1447 ;
        RECT 0.112 0.3673 0.144 0.3887 ;
        RECT 0.112 0.3887 0.144 0.4467 ;
        RECT 0.144 0.1233 0.157 0.1447 ;
        RECT 0.144 0.3673 0.157 0.3887 ;
        RECT 0.144 0.3887 0.157 0.4467 ;
        RECT 0.157 0.1233 0.462 0.1447 ;
        RECT 0.157 0.3673 0.462 0.3887 ;
        RECT 0.462 0.1233 0.49 0.1447 ;
        RECT 0.462 0.1447 0.49 0.2467 ;
        RECT 0.462 0.2467 0.49 0.2653 ;
        RECT 0.462 0.2653 0.49 0.3673 ;
        RECT 0.462 0.3673 0.49 0.3887 ;
        RECT 0.49 0.2467 1.07 0.2653 ;
      LAYER M1 ;
        RECT 0.098 0.3673 0.112 0.3887 ;
        RECT 0.098 0.3887 0.112 0.4467 ;
        RECT 0.112 0.0653 0.144 0.1233 ;
        RECT 0.112 0.1233 0.144 0.1447 ;
        RECT 0.112 0.3673 0.144 0.3887 ;
        RECT 0.112 0.3887 0.144 0.4467 ;
        RECT 0.144 0.1233 0.157 0.1447 ;
        RECT 0.144 0.3673 0.157 0.3887 ;
        RECT 0.144 0.3887 0.157 0.4467 ;
        RECT 0.157 0.1233 0.462 0.1447 ;
        RECT 0.157 0.3673 0.462 0.3887 ;
        RECT 0.462 0.1233 0.49 0.1447 ;
        RECT 0.462 0.1447 0.49 0.2467 ;
        RECT 0.462 0.2467 0.49 0.2653 ;
        RECT 0.462 0.2653 0.49 0.3673 ;
        RECT 0.462 0.3673 0.49 0.3887 ;
        RECT 0.49 0.2467 1.07 0.2653 ;
  END
END BUF_X12_8T

MACRO BUF_X16_8T
  CLASS core ;
  FOREIGN BUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1547 0.078 0.2367 ;
        RECT 0.05 0.2367 0.078 0.2753 ;
        RECT 0.05 0.2753 0.078 0.3413 ;
        RECT 0.078 0.2367 0.554 0.2753 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0679 1.454 0.0867 ;
        RECT 0.594 0.4213 1.454 0.44 ;
        RECT 1.454 0.0679 1.52 0.0867 ;
        RECT 1.454 0.4213 1.52 0.44 ;
        RECT 1.52 0.0679 1.552 0.0867 ;
        RECT 1.52 0.0867 1.552 0.4213 ;
        RECT 1.52 0.4213 1.552 0.44 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.454 0.5307 ;
        RECT 1.454 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0653 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.3053 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.4287 ;
        RECT 0.1419 0.1367 0.59 0.1553 ;
        RECT 0.1419 0.3053 0.59 0.324 ;
        RECT 0.59 0.1367 0.618 0.1553 ;
        RECT 0.59 0.1553 0.618 0.2453 ;
        RECT 0.59 0.2453 0.618 0.264 ;
        RECT 0.59 0.264 0.618 0.3053 ;
        RECT 0.59 0.3053 0.618 0.324 ;
        RECT 0.618 0.2453 1.454 0.264 ;
      LAYER M1 ;
        RECT 0.114 0.0653 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.3053 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.4287 ;
        RECT 0.1419 0.1367 0.59 0.1553 ;
        RECT 0.1419 0.3053 0.59 0.324 ;
        RECT 0.59 0.1367 0.618 0.1553 ;
        RECT 0.59 0.1553 0.618 0.2453 ;
        RECT 0.59 0.2453 0.618 0.264 ;
        RECT 0.59 0.264 0.618 0.3053 ;
        RECT 0.59 0.3053 0.618 0.324 ;
        RECT 0.618 0.2453 1.454 0.264 ;
  END
END BUF_X16_8T

MACRO CLKBUF_X1_8T
  CLASS core ;
  FOREIGN CLKBUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.076 0.272 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1429 0.5307 ;
        RECT 0.1429 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.262 0.115 0.3053 ;
        RECT 0.114 0.3053 0.115 0.3487 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.262 ;
        RECT 0.115 0.262 0.1419 0.3053 ;
        RECT 0.115 0.3053 0.1419 0.3487 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.262 ;
        RECT 0.1419 0.262 0.1429 0.3053 ;
      LAYER M1 ;
        RECT 0.114 0.048 0.115 0.1233 ;
        RECT 0.114 0.1233 0.115 0.142 ;
        RECT 0.114 0.262 0.115 0.3053 ;
        RECT 0.114 0.3053 0.115 0.3487 ;
        RECT 0.115 0.048 0.1419 0.1233 ;
        RECT 0.115 0.1233 0.1419 0.142 ;
        RECT 0.115 0.142 0.1419 0.262 ;
        RECT 0.115 0.262 0.1419 0.3053 ;
        RECT 0.115 0.3053 0.1419 0.3487 ;
        RECT 0.1419 0.1233 0.1429 0.142 ;
        RECT 0.1419 0.142 0.1429 0.262 ;
        RECT 0.1419 0.262 0.1429 0.3053 ;
  END
END CLKBUF_X1_8T

MACRO CLKBUF_X2_8T
  CLASS core ;
  FOREIGN CLKBUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1973 0.078 0.3413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.4253 0.178 0.4693 ;
        RECT 0.178 0.048 0.206 0.4253 ;
        RECT 0.178 0.4253 0.206 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.086 0.08 0.128 ;
        RECT 0.048 0.128 0.08 0.1467 ;
        RECT 0.048 0.3707 0.08 0.3893 ;
        RECT 0.048 0.3893 0.08 0.4573 ;
        RECT 0.08 0.128 0.114 0.1467 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
      LAYER M1 ;
        RECT 0.048 0.086 0.08 0.128 ;
        RECT 0.048 0.128 0.08 0.1467 ;
        RECT 0.048 0.3707 0.08 0.3893 ;
        RECT 0.048 0.3893 0.08 0.4573 ;
        RECT 0.08 0.128 0.114 0.1467 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.128 0.1419 0.1467 ;
        RECT 0.114 0.1467 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
  END
END CLKBUF_X2_8T

MACRO CLKBUF_X4_8T
  CLASS core ;
  FOREIGN CLKBUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3507 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.0679 0.205 0.0867 ;
        RECT 0.205 0.0679 0.206 0.0867 ;
        RECT 0.205 0.4253 0.206 0.444 ;
        RECT 0.206 0.0679 0.368 0.0867 ;
        RECT 0.206 0.4253 0.368 0.444 ;
        RECT 0.368 0.0679 0.4 0.0867 ;
        RECT 0.368 0.0867 0.4 0.4253 ;
        RECT 0.368 0.4253 0.4 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.041 0.1107 0.082 0.1293 ;
        RECT 0.082 0.1107 0.178 0.1293 ;
        RECT 0.082 0.3827 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.3827 ;
        RECT 0.178 0.3827 0.206 0.4013 ;
      LAYER M1 ;
        RECT 0.041 0.1107 0.082 0.1293 ;
        RECT 0.082 0.1107 0.178 0.1293 ;
        RECT 0.082 0.3827 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.3827 ;
        RECT 0.178 0.3827 0.206 0.4013 ;
  END
END CLKBUF_X4_8T

MACRO CLKBUF_X8_8T
  CLASS core ;
  FOREIGN CLKBUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.2187 ;
        RECT 0.05 0.2187 0.078 0.2373 ;
        RECT 0.05 0.2373 0.078 0.3413 ;
        RECT 0.078 0.1707 0.079 0.2187 ;
        RECT 0.078 0.2187 0.079 0.2373 ;
        RECT 0.079 0.2187 0.318 0.2373 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.0679 0.718 0.0867 ;
        RECT 0.338 0.4253 0.718 0.444 ;
        RECT 0.718 0.0679 0.754 0.0867 ;
        RECT 0.718 0.4253 0.754 0.444 ;
        RECT 0.754 0.0679 0.782 0.0867 ;
        RECT 0.754 0.0867 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3 0.1419 0.3213 ;
        RECT 0.114 0.3213 0.1419 0.3613 ;
        RECT 0.1419 0.1107 0.406 0.1293 ;
        RECT 0.1419 0.3 0.406 0.3213 ;
        RECT 0.406 0.1107 0.434 0.1293 ;
        RECT 0.406 0.1293 0.434 0.238 ;
        RECT 0.406 0.238 0.434 0.2767 ;
        RECT 0.406 0.2767 0.434 0.3 ;
        RECT 0.406 0.3 0.434 0.3213 ;
        RECT 0.434 0.238 0.718 0.2767 ;
      LAYER M1 ;
        RECT 0.05 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3 0.1419 0.3213 ;
        RECT 0.114 0.3213 0.1419 0.3613 ;
        RECT 0.1419 0.1107 0.406 0.1293 ;
        RECT 0.1419 0.3 0.406 0.3213 ;
        RECT 0.406 0.1107 0.434 0.1293 ;
        RECT 0.406 0.1293 0.434 0.238 ;
        RECT 0.406 0.238 0.434 0.2767 ;
        RECT 0.406 0.2767 0.434 0.3 ;
        RECT 0.406 0.3 0.434 0.3213 ;
        RECT 0.434 0.238 0.718 0.2767 ;
  END
END CLKBUF_X8_8T

MACRO CLKBUF_X12_8T
  CLASS core ;
  FOREIGN CLKBUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.1587 0.083 0.224 ;
        RECT 0.045 0.224 0.083 0.2453 ;
        RECT 0.045 0.2453 0.083 0.3533 ;
        RECT 0.083 0.224 0.426 0.2453 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.0679 0.998 0.0867 ;
        RECT 0.466 0.4253 0.998 0.444 ;
        RECT 0.998 0.0679 1.1359 0.0867 ;
        RECT 0.998 0.4253 1.1359 0.444 ;
        RECT 1.1359 0.0679 1.168 0.0867 ;
        RECT 1.1359 0.0867 1.168 0.4253 ;
        RECT 1.1359 0.4253 1.168 0.444 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.998 0.5307 ;
        RECT 0.998 0.4933 1.29 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.29 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0429 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3667 0.1419 0.3853 ;
        RECT 0.114 0.3853 0.1419 0.4467 ;
        RECT 0.1419 0.1107 0.462 0.1293 ;
        RECT 0.1419 0.3667 0.462 0.3853 ;
        RECT 0.462 0.1107 0.49 0.1293 ;
        RECT 0.462 0.1293 0.49 0.2093 ;
        RECT 0.462 0.2093 0.49 0.2306 ;
        RECT 0.462 0.2306 0.49 0.3667 ;
        RECT 0.462 0.3667 0.49 0.3853 ;
        RECT 0.49 0.1107 0.494 0.1293 ;
        RECT 0.49 0.1293 0.494 0.2093 ;
        RECT 0.49 0.2093 0.494 0.2306 ;
        RECT 0.494 0.2093 0.998 0.2306 ;
      LAYER M1 ;
        RECT 0.0429 0.1107 0.114 0.1293 ;
        RECT 0.114 0.1107 0.1419 0.1293 ;
        RECT 0.114 0.3667 0.1419 0.3853 ;
        RECT 0.114 0.3853 0.1419 0.4467 ;
        RECT 0.1419 0.1107 0.462 0.1293 ;
        RECT 0.1419 0.3667 0.462 0.3853 ;
        RECT 0.462 0.1107 0.49 0.1293 ;
        RECT 0.462 0.1293 0.49 0.2093 ;
        RECT 0.462 0.2093 0.49 0.2306 ;
        RECT 0.462 0.2306 0.49 0.3667 ;
        RECT 0.462 0.3667 0.49 0.3853 ;
        RECT 0.49 0.1107 0.494 0.1293 ;
        RECT 0.49 0.1293 0.494 0.2093 ;
        RECT 0.49 0.2093 0.494 0.2306 ;
        RECT 0.494 0.2093 0.998 0.2306 ;
  END
END CLKBUF_X12_8T

MACRO CLKBUF_X16_8T
  CLASS core ;
  FOREIGN CLKBUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.148 0.078 0.2173 ;
        RECT 0.05 0.2173 0.078 0.2387 ;
        RECT 0.05 0.2387 0.078 0.3507 ;
        RECT 0.078 0.2173 0.554 0.2387 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0579 1.454 0.0967 ;
        RECT 0.594 0.4153 1.454 0.454 ;
        RECT 1.454 0.0579 1.52 0.0967 ;
        RECT 1.454 0.4153 1.52 0.454 ;
        RECT 1.52 0.0579 1.552 0.0967 ;
        RECT 1.52 0.0967 1.552 0.4153 ;
        RECT 1.52 0.4153 1.552 0.454 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.454 0.5307 ;
        RECT 1.454 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0727 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.35 0.1419 0.3753 ;
        RECT 0.114 0.3753 0.1419 0.4253 ;
        RECT 0.1419 0.1367 0.595 0.1553 ;
        RECT 0.1419 0.35 0.595 0.3753 ;
        RECT 0.595 0.1367 0.653 0.1553 ;
        RECT 0.595 0.1553 0.653 0.2107 ;
        RECT 0.595 0.2107 0.653 0.2293 ;
        RECT 0.595 0.2293 0.653 0.35 ;
        RECT 0.595 0.35 0.653 0.3753 ;
        RECT 0.653 0.2107 1.454 0.2293 ;
      LAYER M1 ;
        RECT 0.114 0.0727 0.1419 0.1367 ;
        RECT 0.114 0.1367 0.1419 0.1553 ;
        RECT 0.114 0.35 0.1419 0.3753 ;
        RECT 0.114 0.3753 0.1419 0.4253 ;
        RECT 0.1419 0.1367 0.595 0.1553 ;
        RECT 0.1419 0.35 0.595 0.3753 ;
        RECT 0.595 0.1367 0.653 0.1553 ;
        RECT 0.595 0.1553 0.653 0.2107 ;
        RECT 0.595 0.2107 0.653 0.2293 ;
        RECT 0.595 0.2293 0.653 0.35 ;
        RECT 0.595 0.35 0.653 0.3753 ;
        RECT 0.653 0.2107 1.454 0.2293 ;
  END
END CLKBUF_X16_8T

MACRO CLKGATETST_X1_8T
  CLASS core ;
  FOREIGN CLKGATETST_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.512 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.1587 0.718 0.3413 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.448 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.2133 0.078 0.448 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.01 0.064 1.038 0.436 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.366 0.5307 ;
        RECT 0.366 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.098 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.098 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.21 0.268 0.686 0.2867 ;
        RECT 0.146 0.3107 0.522 0.3293 ;
        RECT 0.73 0.268 1.006 0.2867 ;
      LAYER MINT1 ;
        RECT 0.21 0.268 0.686 0.2867 ;
        RECT 0.146 0.3107 0.522 0.3293 ;
        RECT 0.73 0.268 1.006 0.2867 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.238 0.0867 ;
        RECT 0.242 0.176 0.27 0.3607 ;
        RECT 0.37 0.1613 0.398 0.3347 ;
        RECT 0.462 0.248 0.494 0.34 ;
        RECT 0.626 0.1107 0.654 0.1293 ;
        RECT 0.626 0.1293 0.654 0.3707 ;
        RECT 0.626 0.3707 0.654 0.3947 ;
        RECT 0.654 0.1107 0.75 0.1293 ;
        RECT 0.654 0.3707 0.75 0.3947 ;
        RECT 0.75 0.1107 0.755 0.1293 ;
        RECT 0.754 0.1653 0.79 0.3087 ;
        RECT 0.754 0.3087 0.79 0.3347 ;
        RECT 0.79 0.3087 0.8179 0.3347 ;
        RECT 0.8179 0.3087 0.846 0.3347 ;
        RECT 0.8179 0.3347 0.846 0.3893 ;
        RECT 0.946 0.1507 0.974 0.3827 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.4187 ;
        RECT 0.178 0.4187 0.206 0.4507 ;
        RECT 0.206 0.1107 0.302 0.1293 ;
        RECT 0.206 0.4187 0.302 0.4507 ;
        RECT 0.302 0.4187 0.366 0.4507 ;
        RECT 0.306 0.2047 0.334 0.364 ;
        RECT 0.306 0.364 0.334 0.3827 ;
        RECT 0.334 0.364 0.558 0.3827 ;
        RECT 0.558 0.1227 0.59 0.2047 ;
        RECT 0.558 0.2047 0.59 0.364 ;
        RECT 0.558 0.364 0.59 0.3827 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.2227 ;
        RECT 0.462 0.0679 0.466 0.0867 ;
        RECT 0.466 0.0679 0.882 0.0867 ;
        RECT 0.466 0.4187 0.882 0.4507 ;
        RECT 0.882 0.0679 0.91 0.0867 ;
        RECT 0.882 0.0867 0.91 0.2227 ;
        RECT 0.882 0.2227 0.91 0.4187 ;
        RECT 0.882 0.4187 0.91 0.4507 ;
      LAYER V1 ;
        RECT 0.178 0.3107 0.206 0.3293 ;
        RECT 0.242 0.268 0.27 0.2867 ;
        RECT 0.37 0.268 0.398 0.2867 ;
        RECT 0.462 0.3107 0.49 0.3293 ;
        RECT 0.626 0.268 0.654 0.2867 ;
        RECT 0.762 0.268 0.79 0.2867 ;
        RECT 0.946 0.268 0.974 0.2867 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.238 0.0867 ;
        RECT 0.242 0.176 0.27 0.3607 ;
        RECT 0.37 0.1613 0.398 0.3347 ;
        RECT 0.462 0.248 0.494 0.34 ;
        RECT 0.626 0.1107 0.654 0.1293 ;
        RECT 0.626 0.1293 0.654 0.3707 ;
        RECT 0.626 0.3707 0.654 0.3947 ;
        RECT 0.654 0.1107 0.75 0.1293 ;
        RECT 0.654 0.3707 0.75 0.3947 ;
        RECT 0.75 0.1107 0.755 0.1293 ;
        RECT 0.754 0.1653 0.79 0.3087 ;
        RECT 0.754 0.3087 0.79 0.3347 ;
        RECT 0.79 0.3087 0.8179 0.3347 ;
        RECT 0.8179 0.3087 0.846 0.3347 ;
        RECT 0.8179 0.3347 0.846 0.3893 ;
        RECT 0.946 0.1507 0.974 0.3827 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.4187 ;
        RECT 0.178 0.4187 0.206 0.4507 ;
        RECT 0.206 0.1107 0.302 0.1293 ;
        RECT 0.206 0.4187 0.302 0.4507 ;
        RECT 0.302 0.4187 0.366 0.4507 ;
        RECT 0.306 0.2047 0.334 0.364 ;
        RECT 0.306 0.364 0.334 0.3827 ;
        RECT 0.334 0.364 0.558 0.3827 ;
        RECT 0.558 0.1227 0.59 0.2047 ;
        RECT 0.558 0.2047 0.59 0.364 ;
        RECT 0.558 0.364 0.59 0.3827 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.2227 ;
        RECT 0.462 0.0679 0.466 0.0867 ;
        RECT 0.466 0.0679 0.882 0.0867 ;
        RECT 0.466 0.4187 0.882 0.4507 ;
        RECT 0.882 0.0679 0.91 0.0867 ;
        RECT 0.882 0.0867 0.91 0.2227 ;
        RECT 0.882 0.2227 0.91 0.4187 ;
        RECT 0.882 0.4187 0.91 0.4507 ;
  END
END CLKGATETST_X1_8T

MACRO DFFRNQ_X1_8T
  CLASS core ;
  FOREIGN DFFRNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.1827 1.1339 0.2013 ;
        RECT 1.1339 0.1827 1.326 0.2013 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.0427 1.616 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.8139 0.5307 ;
        RECT 0.8139 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.102 0.5307 ;
        RECT 1.102 0.4933 1.188 0.5307 ;
        RECT 1.188 0.4933 1.488 0.5307 ;
        RECT 1.488 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.53 0.4153 0.8139 0.454 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.292 ;
        RECT 0.434 0.292 0.462 0.4467 ;
        RECT 0.462 0.0679 0.8 0.0867 ;
        RECT 0.8 0.0679 0.828 0.0867 ;
        RECT 0.8 0.0867 0.828 0.292 ;
        RECT 0.576 0.22 0.604 0.3373 ;
        RECT 0.576 0.3373 0.604 0.356 ;
        RECT 0.604 0.3373 0.882 0.356 ;
        RECT 0.882 0.048 0.91 0.22 ;
        RECT 0.882 0.22 0.91 0.3373 ;
        RECT 0.882 0.3373 0.91 0.356 ;
        RECT 0.882 0.356 0.91 0.448 ;
        RECT 1.01 0.0679 1.038 0.0867 ;
        RECT 1.01 0.0867 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.4467 ;
        RECT 1.038 0.0679 1.335 0.0867 ;
        RECT 1.335 0.0679 1.363 0.0867 ;
        RECT 1.335 0.0867 1.363 0.244 ;
        RECT 1.224 0.2627 1.252 0.4253 ;
        RECT 1.224 0.4253 1.252 0.444 ;
        RECT 1.252 0.4253 1.458 0.444 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.4253 ;
        RECT 1.458 0.4253 1.486 0.444 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.4253 ;
        RECT 1.486 0.4253 1.488 0.444 ;
        RECT 0.048 0.0567 0.08 0.0939 ;
        RECT 0.048 0.0939 0.08 0.1127 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0939 0.114 0.1127 ;
        RECT 0.08 0.3779 0.114 0.404 ;
        RECT 0.114 0.0939 0.1419 0.1127 ;
        RECT 0.114 0.1127 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3827 ;
        RECT 0.526 0.1293 0.558 0.196 ;
        RECT 0.736 0.172 0.764 0.292 ;
        RECT 0.946 0.1827 0.974 0.3853 ;
        RECT 1.074 0.1159 1.102 0.2113 ;
        RECT 1.074 0.3067 1.102 0.4147 ;
        RECT 1.156 0.1107 1.188 0.4573 ;
        RECT 1.266 0.1159 1.294 0.212 ;
      LAYER V1 ;
        RECT 0.114 0.3533 0.1419 0.372 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.37 0.14 0.398 0.1587 ;
        RECT 0.498 0.3533 0.526 0.372 ;
        RECT 0.53 0.14 0.558 0.1587 ;
        RECT 0.736 0.1827 0.764 0.2013 ;
        RECT 0.946 0.3533 0.974 0.372 ;
        RECT 1.074 0.14 1.102 0.1587 ;
        RECT 1.074 0.3533 1.102 0.372 ;
        RECT 1.266 0.1827 1.294 0.2013 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.53 0.4153 0.8139 0.454 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.292 ;
        RECT 0.434 0.292 0.462 0.4467 ;
        RECT 0.462 0.0679 0.8 0.0867 ;
        RECT 0.8 0.0679 0.828 0.0867 ;
        RECT 0.8 0.0867 0.828 0.292 ;
        RECT 0.576 0.22 0.604 0.3373 ;
        RECT 0.576 0.3373 0.604 0.356 ;
        RECT 0.604 0.3373 0.882 0.356 ;
        RECT 0.882 0.048 0.91 0.22 ;
        RECT 0.882 0.22 0.91 0.3373 ;
        RECT 0.882 0.3373 0.91 0.356 ;
        RECT 0.882 0.356 0.91 0.448 ;
        RECT 1.01 0.0679 1.038 0.0867 ;
        RECT 1.01 0.0867 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.4467 ;
        RECT 1.038 0.0679 1.335 0.0867 ;
        RECT 1.335 0.0679 1.363 0.0867 ;
        RECT 1.335 0.0867 1.363 0.244 ;
        RECT 1.224 0.2627 1.252 0.4253 ;
        RECT 1.224 0.4253 1.252 0.444 ;
        RECT 1.252 0.4253 1.458 0.444 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.4253 ;
        RECT 1.458 0.4253 1.486 0.444 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.4253 ;
        RECT 1.486 0.4253 1.488 0.444 ;
        RECT 0.048 0.0567 0.08 0.0939 ;
        RECT 0.048 0.0939 0.08 0.1127 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0939 0.114 0.1127 ;
        RECT 0.08 0.3779 0.114 0.404 ;
        RECT 0.114 0.0939 0.1419 0.1127 ;
        RECT 0.114 0.1127 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3827 ;
        RECT 0.526 0.1293 0.558 0.196 ;
        RECT 0.736 0.172 0.764 0.292 ;
        RECT 0.946 0.1827 0.974 0.3853 ;
        RECT 1.074 0.1159 1.102 0.2113 ;
        RECT 1.074 0.3067 1.102 0.4147 ;
        RECT 1.156 0.1107 1.188 0.4573 ;
        RECT 1.266 0.1159 1.294 0.212 ;
  END
END DFFRNQ_X1_8T

MACRO DFFSNQ_X1_8T
  CLASS core ;
  FOREIGN DFFSNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.1827 1.1339 0.2013 ;
        RECT 1.1339 0.1827 1.326 0.2013 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.0427 1.616 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.554 0.5307 ;
        RECT 0.554 0.4933 0.91 0.5307 ;
        RECT 0.91 0.4933 0.974 0.5307 ;
        RECT 0.974 0.4933 1.106 0.5307 ;
        RECT 1.106 0.4933 1.3899 0.5307 ;
        RECT 1.3899 0.4933 1.488 0.5307 ;
        RECT 1.488 0.4933 1.674 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.674 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER MINT1 ;
        RECT 0.146 0.14 1.1339 0.1587 ;
        RECT 0.082 0.3533 1.1339 0.372 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.434 0.0813 0.462 0.1 ;
        RECT 0.434 0.1 0.462 0.244 ;
        RECT 0.434 0.244 0.462 0.4467 ;
        RECT 0.462 0.0813 0.8179 0.1 ;
        RECT 0.8179 0.0813 0.846 0.1 ;
        RECT 0.8179 0.1 0.846 0.244 ;
        RECT 0.946 0.1827 0.974 0.3827 ;
        RECT 1.074 0.1293 1.106 0.2167 ;
        RECT 1.074 0.262 1.106 0.396 ;
        RECT 1.266 0.124 1.294 0.212 ;
        RECT 1.202 0.2627 1.23 0.3827 ;
        RECT 1.202 0.3827 1.23 0.4013 ;
        RECT 1.23 0.3827 1.458 0.4013 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.3827 ;
        RECT 1.458 0.3827 1.486 0.4013 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.3827 ;
        RECT 1.486 0.3827 1.488 0.4013 ;
        RECT 0.045 0.0547 0.048 0.092 ;
        RECT 0.045 0.092 0.048 0.118 ;
        RECT 0.048 0.0547 0.08 0.092 ;
        RECT 0.048 0.092 0.08 0.118 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0547 0.083 0.092 ;
        RECT 0.08 0.092 0.083 0.118 ;
        RECT 0.08 0.3779 0.083 0.404 ;
        RECT 0.083 0.092 0.114 0.118 ;
        RECT 0.083 0.3779 0.114 0.404 ;
        RECT 0.114 0.092 0.1419 0.118 ;
        RECT 0.114 0.118 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3933 ;
        RECT 0.526 0.1293 0.554 0.2033 ;
        RECT 0.754 0.172 0.782 0.244 ;
        RECT 0.608 0.1827 0.636 0.3827 ;
        RECT 0.608 0.3827 0.636 0.4013 ;
        RECT 0.636 0.3827 0.878 0.4013 ;
        RECT 0.878 0.3827 0.882 0.4013 ;
        RECT 0.878 0.4013 0.882 0.4573 ;
        RECT 0.882 0.064 0.91 0.1827 ;
        RECT 0.882 0.1827 0.91 0.3827 ;
        RECT 0.882 0.3827 0.91 0.4013 ;
        RECT 0.882 0.4013 0.91 0.4573 ;
        RECT 1.01 0.076 1.038 0.0946 ;
        RECT 1.01 0.0946 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.448 ;
        RECT 1.038 0.076 1.352 0.0946 ;
        RECT 1.352 0.076 1.3799 0.0946 ;
        RECT 1.352 0.0946 1.3799 0.244 ;
        RECT 1.106 0.4253 1.3899 0.444 ;
      LAYER V1 ;
        RECT 0.114 0.3533 0.1419 0.372 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.37 0.14 0.398 0.1587 ;
        RECT 0.498 0.3533 0.526 0.372 ;
        RECT 0.526 0.14 0.554 0.1587 ;
        RECT 0.754 0.1827 0.782 0.2013 ;
        RECT 0.946 0.3533 0.974 0.372 ;
        RECT 1.074 0.14 1.102 0.1587 ;
        RECT 1.074 0.3533 1.102 0.372 ;
        RECT 1.266 0.1827 1.294 0.2013 ;
      LAYER M1 ;
        RECT 0.178 0.048 0.206 0.4639 ;
        RECT 0.306 0.048 0.334 0.4639 ;
        RECT 0.434 0.0813 0.462 0.1 ;
        RECT 0.434 0.1 0.462 0.244 ;
        RECT 0.434 0.244 0.462 0.4467 ;
        RECT 0.462 0.0813 0.8179 0.1 ;
        RECT 0.8179 0.0813 0.846 0.1 ;
        RECT 0.8179 0.1 0.846 0.244 ;
        RECT 0.946 0.1827 0.974 0.3827 ;
        RECT 1.074 0.1293 1.106 0.2167 ;
        RECT 1.074 0.262 1.106 0.396 ;
        RECT 1.266 0.124 1.294 0.212 ;
        RECT 1.202 0.2627 1.23 0.3827 ;
        RECT 1.202 0.3827 1.23 0.4013 ;
        RECT 1.23 0.3827 1.458 0.4013 ;
        RECT 1.458 0.048 1.486 0.088 ;
        RECT 1.458 0.088 1.486 0.2627 ;
        RECT 1.458 0.2627 1.486 0.3827 ;
        RECT 1.458 0.3827 1.486 0.4013 ;
        RECT 1.486 0.088 1.488 0.2627 ;
        RECT 1.486 0.2627 1.488 0.3827 ;
        RECT 1.486 0.3827 1.488 0.4013 ;
        RECT 0.045 0.0547 0.048 0.092 ;
        RECT 0.045 0.092 0.048 0.118 ;
        RECT 0.048 0.0547 0.08 0.092 ;
        RECT 0.048 0.092 0.08 0.118 ;
        RECT 0.048 0.3779 0.08 0.404 ;
        RECT 0.048 0.404 0.08 0.4573 ;
        RECT 0.08 0.0547 0.083 0.092 ;
        RECT 0.08 0.092 0.083 0.118 ;
        RECT 0.08 0.3779 0.083 0.404 ;
        RECT 0.083 0.092 0.114 0.118 ;
        RECT 0.083 0.3779 0.114 0.404 ;
        RECT 0.114 0.092 0.1419 0.118 ;
        RECT 0.114 0.118 0.1419 0.3779 ;
        RECT 0.114 0.3779 0.1419 0.404 ;
        RECT 0.37 0.1293 0.398 0.3293 ;
        RECT 0.498 0.268 0.526 0.3933 ;
        RECT 0.526 0.1293 0.554 0.2033 ;
        RECT 0.754 0.172 0.782 0.244 ;
        RECT 0.608 0.1827 0.636 0.3827 ;
        RECT 0.608 0.3827 0.636 0.4013 ;
        RECT 0.636 0.3827 0.878 0.4013 ;
        RECT 0.878 0.3827 0.882 0.4013 ;
        RECT 0.878 0.4013 0.882 0.4573 ;
        RECT 0.882 0.064 0.91 0.1827 ;
        RECT 0.882 0.1827 0.91 0.3827 ;
        RECT 0.882 0.3827 0.91 0.4013 ;
        RECT 0.882 0.4013 0.91 0.4573 ;
        RECT 1.01 0.076 1.038 0.0946 ;
        RECT 1.01 0.0946 1.038 0.244 ;
        RECT 1.01 0.244 1.038 0.448 ;
        RECT 1.038 0.076 1.352 0.0946 ;
        RECT 1.352 0.076 1.3799 0.0946 ;
        RECT 1.352 0.0946 1.3799 0.244 ;
        RECT 1.106 0.4253 1.3899 0.444 ;
  END
END DFFSNQ_X1_8T

MACRO FA_X1_8T
  CLASS core ;
  FOREIGN FA_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.536 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.21 0.3107 1.098 0.3293 ;
      LAYER V1 ;
        RECT 0.656 0.3107 0.684 0.3293 ;
        RECT 1.038 0.3107 1.066 0.3293 ;
      LAYER M1 ;
        RECT 0.656 0.268 0.684 0.3507 ;
        RECT 1.038 0.1827 1.074 0.3507 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.1827 0.1827 0.789 0.2013 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.146 0.14 1.262 0.1587 ;
      LAYER V1 ;
        RECT 0.178 0.14 0.206 0.1587 ;
        RECT 0.58 0.14 0.608 0.1587 ;
        RECT 1.202 0.14 1.23 0.1587 ;
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3933 ;
        RECT 0.58 0.1293 0.608 0.244 ;
        RECT 1.202 0.1187 1.23 0.244 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.458 0.076 1.486 0.436 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.138 0.846 0.4267 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.767 0.5307 ;
        RECT 0.767 0.4933 1.038 0.5307 ;
        RECT 1.038 0.4933 1.084 0.5307 ;
        RECT 1.084 0.4933 1.166 0.5307 ;
        RECT 1.166 0.4933 1.289 0.5307 ;
        RECT 1.289 0.4933 1.358 0.5307 ;
        RECT 1.358 0.4933 1.546 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.546 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.082 0.268 1.321 0.2867 ;
        RECT 0.402 0.2253 1.3899 0.244 ;
      LAYER MINT1 ;
        RECT 0.082 0.268 1.321 0.2867 ;
        RECT 0.402 0.2253 1.3899 0.244 ;
      LAYER M1 ;
        RECT 0.027 0.1187 0.065 0.2253 ;
        RECT 0.027 0.2253 0.065 0.244 ;
        RECT 0.065 0.2253 0.103 0.244 ;
        RECT 0.103 0.2253 0.1419 0.244 ;
        RECT 0.103 0.244 0.1419 0.308 ;
        RECT 0.242 0.1827 0.27 0.3933 ;
        RECT 0.424 0.1827 0.462 0.338 ;
        RECT 0.37 0.0647 0.618 0.09 ;
        RECT 0.37 0.3833 0.402 0.402 ;
        RECT 0.37 0.402 0.402 0.4653 ;
        RECT 0.402 0.3833 0.624 0.402 ;
        RECT 0.624 0.3833 0.656 0.402 ;
        RECT 0.624 0.402 0.656 0.4653 ;
        RECT 0.624 0.4653 0.656 0.4693 ;
        RECT 0.729 0.1627 0.767 0.3093 ;
        RECT 0.882 0.1293 0.91 0.244 ;
        RECT 0.882 0.3747 0.91 0.3933 ;
        RECT 0.882 0.3933 0.91 0.4639 ;
        RECT 0.91 0.3747 1.01 0.3933 ;
        RECT 1.01 0.3747 1.038 0.3933 ;
        RECT 1.01 0.3933 1.038 0.4639 ;
        RECT 1.1379 0.048 1.166 0.4639 ;
        RECT 1.2609 0.2573 1.289 0.3933 ;
        RECT 0.306 0.064 0.334 0.448 ;
        RECT 0.498 0.1827 0.526 0.338 ;
        RECT 0.946 0.1827 0.984 0.3293 ;
        RECT 0.846 0.0667 1.084 0.066732 ;
        RECT 1.33 0.1827 1.358 0.3507 ;
      LAYER V1 ;
        RECT 0.114 0.268 0.1419 0.2867 ;
        RECT 0.242 0.3107 0.27 0.3293 ;
        RECT 0.306 0.1827 0.334 0.2013 ;
        RECT 0.434 0.2253 0.462 0.244 ;
        RECT 0.498 0.268 0.526 0.2867 ;
        RECT 0.729 0.1827 0.757 0.2013 ;
        RECT 0.882 0.14 0.91 0.1587 ;
        RECT 0.956 0.268 0.984 0.2867 ;
        RECT 1.1379 0.2253 1.166 0.244 ;
        RECT 1.2609 0.268 1.289 0.2867 ;
        RECT 1.33 0.2253 1.358 0.244 ;
      LAYER M1 ;
        RECT 0.027 0.1187 0.065 0.2253 ;
        RECT 0.027 0.2253 0.065 0.244 ;
        RECT 0.065 0.2253 0.103 0.244 ;
        RECT 0.103 0.2253 0.1419 0.244 ;
        RECT 0.103 0.244 0.1419 0.308 ;
        RECT 0.242 0.1827 0.27 0.3933 ;
        RECT 0.424 0.1827 0.462 0.338 ;
        RECT 0.37 0.0647 0.618 0.09 ;
        RECT 0.37 0.3833 0.402 0.402 ;
        RECT 0.37 0.402 0.402 0.4653 ;
        RECT 0.402 0.3833 0.624 0.402 ;
        RECT 0.624 0.3833 0.656 0.402 ;
        RECT 0.624 0.402 0.656 0.4653 ;
        RECT 0.624 0.4653 0.656 0.4693 ;
        RECT 0.729 0.1627 0.767 0.3093 ;
        RECT 0.882 0.1293 0.91 0.244 ;
        RECT 0.882 0.3747 0.91 0.3933 ;
        RECT 0.882 0.3933 0.91 0.4639 ;
        RECT 0.91 0.3747 1.01 0.3933 ;
        RECT 1.01 0.3747 1.038 0.3933 ;
        RECT 1.01 0.3933 1.038 0.4639 ;
        RECT 1.1379 0.048 1.166 0.4639 ;
        RECT 1.2609 0.2573 1.289 0.3933 ;
        RECT 0.306 0.064 0.334 0.448 ;
        RECT 0.498 0.1827 0.526 0.338 ;
        RECT 0.946 0.1827 0.984 0.3293 ;
        RECT 0.846 0.0667 1.084 0.066732 ;
        RECT 1.33 0.1827 1.358 0.3507 ;
  END
END FA_X1_8T

MACRO FILLTIE_8T
  CLASS core ;
  FOREIGN FILLTIE_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.578 BY 0.512 ;
  OBS
      LAYER M1 ;
        RECT -0.01 -0.0187 0.588 0.0187 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
      LAYER M1 ;
        RECT -0.01 -0.0187 0.588 0.0187 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
  END
END FILLTIE_8T

MACRO FILL_X1_8T
  CLASS core ;
  FOREIGN FILL_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.128 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.138 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.138 0.0187 ;
    END
  END VSS
END FILL_X1_8T

MACRO FILL_X2_8T
  CLASS core ;
  FOREIGN FILL_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
END FILL_X2_8T

MACRO FILL_X4_8T
  CLASS core ;
  FOREIGN FILL_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.33 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.33 0.0187 ;
    END
  END VSS
END FILL_X4_8T

MACRO FILL_X8_8T
  CLASS core ;
  FOREIGN FILL_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
END FILL_X8_8T

MACRO FILL_X16_8T
  CLASS core ;
  FOREIGN FILL_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.512 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.098 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.098 0.0187 ;
    END
  END VSS
END FILL_X16_8T

MACRO HA_X1_8T
  CLASS core ;
  FOREIGN HA_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.512 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1827 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
        RECT 0.27 0.3707 0.434 0.3893 ;
        RECT 0.434 0.1827 0.462 0.3707 ;
        RECT 0.434 0.3707 0.462 0.3893 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.3413 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0547 0.078 0.4253 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.754 0.12 0.782 0.4253 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.596 0.5307 ;
        RECT 0.596 0.4933 0.66 0.5307 ;
        RECT 0.66 0.4933 0.842 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.842 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.338 0.0679 0.622 0.0867 ;
        RECT 0.406 0.1227 0.498 0.144 ;
        RECT 0.498 0.1227 0.53 0.144 ;
        RECT 0.498 0.144 0.53 0.308 ;
        RECT 0.498 0.308 0.53 0.4013 ;
        RECT 0.53 0.1227 0.632 0.144 ;
        RECT 0.632 0.1227 0.66 0.144 ;
        RECT 0.632 0.144 0.66 0.308 ;
        RECT 0.114 0.1107 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.1827 ;
        RECT 0.114 0.1827 0.1419 0.4253 ;
        RECT 0.114 0.4253 0.1419 0.444 ;
        RECT 0.1419 0.1107 0.37 0.132 ;
        RECT 0.1419 0.4253 0.37 0.444 ;
        RECT 0.37 0.4253 0.5659 0.444 ;
        RECT 0.5659 0.1827 0.596 0.4253 ;
        RECT 0.5659 0.4253 0.596 0.444 ;
      LAYER M1 ;
        RECT 0.338 0.0679 0.622 0.0867 ;
        RECT 0.406 0.1227 0.498 0.144 ;
        RECT 0.498 0.1227 0.53 0.144 ;
        RECT 0.498 0.144 0.53 0.308 ;
        RECT 0.498 0.308 0.53 0.4013 ;
        RECT 0.53 0.1227 0.632 0.144 ;
        RECT 0.632 0.1227 0.66 0.144 ;
        RECT 0.632 0.144 0.66 0.308 ;
        RECT 0.114 0.1107 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.1827 ;
        RECT 0.114 0.1827 0.1419 0.4253 ;
        RECT 0.114 0.4253 0.1419 0.444 ;
        RECT 0.1419 0.1107 0.37 0.132 ;
        RECT 0.1419 0.4253 0.37 0.444 ;
        RECT 0.37 0.4253 0.5659 0.444 ;
        RECT 0.5659 0.1827 0.596 0.4253 ;
        RECT 0.5659 0.4253 0.596 0.444 ;
  END
END HA_X1_8T

MACRO INV_X1_8T
  CLASS core ;
  FOREIGN INV_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.076 0.076 0.1419 0.4267 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
END INV_X1_8T

MACRO INV_X2_8T
  CLASS core ;
  FOREIGN INV_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.384 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END INV_X2_8T

MACRO INV_X4_8T
  CLASS core ;
  FOREIGN INV_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.1707 0.08 0.2453 ;
        RECT 0.048 0.2453 0.08 0.264 ;
        RECT 0.048 0.264 0.08 0.3413 ;
        RECT 0.08 0.2453 0.238 0.264 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.0946 0.059 0.1333 ;
        RECT 0.059 0.0946 0.306 0.1333 ;
        RECT 0.059 0.3786 0.306 0.4173 ;
        RECT 0.306 0.0946 0.334 0.1333 ;
        RECT 0.306 0.1333 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4173 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END INV_X4_8T

MACRO INV_X8_8T
  CLASS core ;
  FOREIGN INV_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1293 0.1419 0.264 ;
        RECT 0.114 0.264 0.1419 0.3033 ;
        RECT 0.114 0.3033 0.1419 0.384 ;
        RECT 0.1419 0.264 0.462 0.3033 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.4207 0.054 0.4393 ;
        RECT 0.054 0.0733 0.557 0.092 ;
        RECT 0.054 0.4207 0.557 0.4393 ;
        RECT 0.557 0.0733 0.595 0.092 ;
        RECT 0.557 0.092 0.595 0.4207 ;
        RECT 0.557 0.4207 0.595 0.4393 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
END INV_X8_8T

MACRO INV_X12_8T
  CLASS core ;
  FOREIGN INV_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.2453 ;
        RECT 0.114 0.2453 0.1419 0.264 ;
        RECT 0.114 0.264 0.1419 0.384 ;
        RECT 0.1419 0.2453 0.686 0.264 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.0679 0.8129 0.0867 ;
        RECT 0.054 0.424 0.8129 0.4453 ;
        RECT 0.8129 0.0679 0.851 0.0867 ;
        RECT 0.8129 0.0867 0.851 0.424 ;
        RECT 0.8129 0.424 0.851 0.4453 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
END INV_X12_8T

MACRO LHQ_X1_8T
  CLASS core ;
  FOREIGN LHQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1067 0.27 0.3413 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.0867 0.846 0.4253 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.906 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.906 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.3707 0.05 0.3893 ;
        RECT 0.048 0.3893 0.05 0.4693 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.1227 ;
        RECT 0.05 0.1227 0.078 0.1413 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4693 ;
        RECT 0.078 0.0427 0.08 0.0613 ;
        RECT 0.078 0.1227 0.08 0.1413 ;
        RECT 0.078 0.3707 0.08 0.3893 ;
        RECT 0.078 0.3893 0.08 0.4693 ;
        RECT 0.08 0.0427 0.114 0.0613 ;
        RECT 0.08 0.1227 0.114 0.1413 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.1227 0.1419 0.1413 ;
        RECT 0.114 0.1413 0.1419 0.2147 ;
        RECT 0.114 0.2147 0.1419 0.2333 ;
        RECT 0.114 0.2333 0.1419 0.276 ;
        RECT 0.114 0.276 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0427 0.324 0.0613 ;
        RECT 0.324 0.0427 0.352 0.0613 ;
        RECT 0.324 0.0613 0.352 0.1227 ;
        RECT 0.324 0.1227 0.352 0.1413 ;
        RECT 0.324 0.1413 0.352 0.2147 ;
        RECT 0.324 0.2147 0.23332 0.2333 ;
        RECT 0.23332 0.2147 0.37 0.2333 ;
        RECT 0.37 0.2147 0.398 0.2333 ;
        RECT 0.37 0.2333 0.398 0.276 ;
        RECT 0.53 0.076 0.558 0.0946 ;
        RECT 0.53 0.0946 0.558 0.3293 ;
        RECT 0.558 0.076 0.6899 0.0946 ;
        RECT 0.6899 0.076 0.718 0.0946 ;
        RECT 0.6899 0.0946 0.718 0.3293 ;
        RECT 0.6899 0.3293 0.718 0.3953 ;
        RECT 0.178 0.0907 0.206 0.3067 ;
        RECT 0.178 0.3067 0.206 0.3707 ;
        RECT 0.178 0.3707 0.206 0.3893 ;
        RECT 0.206 0.3707 0.306 0.3893 ;
        RECT 0.306 0.3067 0.34 0.3707 ;
        RECT 0.306 0.3707 0.34 0.3893 ;
        RECT 0.274 0.4253 0.388 0.444 ;
        RECT 0.388 0.076 0.466 0.1153 ;
        RECT 0.388 0.4253 0.466 0.444 ;
        RECT 0.466 0.076 0.494 0.1153 ;
        RECT 0.466 0.1153 0.494 0.204 ;
        RECT 0.466 0.204 0.494 0.4247 ;
        RECT 0.466 0.4247 0.494 0.4253 ;
        RECT 0.466 0.4253 0.494 0.444 ;
        RECT 0.494 0.4247 0.754 0.4253 ;
        RECT 0.494 0.4253 0.754 0.444 ;
        RECT 0.754 0.204 0.782 0.4247 ;
        RECT 0.754 0.4247 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
      LAYER M1 ;
        RECT 0.048 0.3707 0.05 0.3893 ;
        RECT 0.048 0.3893 0.05 0.4693 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.1227 ;
        RECT 0.05 0.1227 0.078 0.1413 ;
        RECT 0.05 0.3707 0.078 0.3893 ;
        RECT 0.05 0.3893 0.078 0.4693 ;
        RECT 0.078 0.0427 0.08 0.0613 ;
        RECT 0.078 0.1227 0.08 0.1413 ;
        RECT 0.078 0.3707 0.08 0.3893 ;
        RECT 0.078 0.3893 0.08 0.4693 ;
        RECT 0.08 0.0427 0.114 0.0613 ;
        RECT 0.08 0.1227 0.114 0.1413 ;
        RECT 0.08 0.3707 0.114 0.3893 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.1227 0.1419 0.1413 ;
        RECT 0.114 0.1413 0.1419 0.2147 ;
        RECT 0.114 0.2147 0.1419 0.2333 ;
        RECT 0.114 0.2333 0.1419 0.276 ;
        RECT 0.114 0.276 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0427 0.324 0.0613 ;
        RECT 0.324 0.0427 0.352 0.0613 ;
        RECT 0.324 0.0613 0.352 0.1227 ;
        RECT 0.324 0.1227 0.352 0.1413 ;
        RECT 0.324 0.1413 0.352 0.2147 ;
        RECT 0.324 0.2147 0.23332 0.2333 ;
        RECT 0.23332 0.2147 0.37 0.2333 ;
        RECT 0.37 0.2147 0.398 0.2333 ;
        RECT 0.37 0.2333 0.398 0.276 ;
        RECT 0.53 0.076 0.558 0.0946 ;
        RECT 0.53 0.0946 0.558 0.3293 ;
        RECT 0.558 0.076 0.6899 0.0946 ;
        RECT 0.6899 0.076 0.718 0.0946 ;
        RECT 0.6899 0.0946 0.718 0.3293 ;
        RECT 0.6899 0.3293 0.718 0.3953 ;
        RECT 0.178 0.0907 0.206 0.3067 ;
        RECT 0.178 0.3067 0.206 0.3707 ;
        RECT 0.178 0.3707 0.206 0.3893 ;
        RECT 0.206 0.3707 0.306 0.3893 ;
        RECT 0.306 0.3067 0.34 0.3707 ;
        RECT 0.306 0.3707 0.34 0.3893 ;
        RECT 0.274 0.4253 0.388 0.444 ;
        RECT 0.388 0.076 0.466 0.1153 ;
        RECT 0.388 0.4253 0.466 0.444 ;
        RECT 0.466 0.076 0.494 0.1153 ;
        RECT 0.466 0.1153 0.494 0.204 ;
        RECT 0.466 0.204 0.494 0.4247 ;
        RECT 0.466 0.4247 0.494 0.4253 ;
        RECT 0.466 0.4253 0.494 0.444 ;
        RECT 0.494 0.4247 0.754 0.4253 ;
        RECT 0.494 0.4253 0.754 0.444 ;
        RECT 0.754 0.204 0.782 0.4247 ;
        RECT 0.754 0.4247 0.782 0.4253 ;
        RECT 0.754 0.4253 0.782 0.444 ;
  END
END LHQ_X1_8T

MACRO MUX2_X1_8T
  CLASS core ;
  FOREIGN MUX2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.512 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.1613 0.59 0.3507 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.2987 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.118 0.4387 0.394 0.4573 ;
      LAYER V1 ;
        RECT 0.15 0.4387 0.206 0.4573 ;
      LAYER M1 ;
        RECT 0.027 0.1613 0.055 0.4387 ;
        RECT 0.027 0.4387 0.055 0.4573 ;
        RECT 0.055 0.4387 0.222 0.4573 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.128 0.718 0.4253 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.842 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.842 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.274 0.2253 0.558 0.244 ;
      LAYER MINT1 ;
        RECT 0.274 0.2253 0.558 0.244 ;
      LAYER M1 ;
        RECT 0.08 0.108 0.099 0.1267 ;
        RECT 0.099 0.108 0.157 0.1267 ;
        RECT 0.099 0.328 0.157 0.3467 ;
        RECT 0.099 0.3467 0.157 0.384 ;
        RECT 0.157 0.108 0.306 0.1267 ;
        RECT 0.157 0.328 0.306 0.3467 ;
        RECT 0.306 0.108 0.334 0.1267 ;
        RECT 0.306 0.1267 0.334 0.328 ;
        RECT 0.306 0.328 0.334 0.3467 ;
        RECT 0.29 0.4387 0.434 0.4693 ;
        RECT 0.434 0.204 0.462 0.4387 ;
        RECT 0.434 0.4387 0.462 0.4693 ;
        RECT 0.498 0.1827 0.526 0.2853 ;
        RECT 0.37 0.0579 0.398 0.0973 ;
        RECT 0.37 0.0973 0.398 0.3293 ;
        RECT 0.37 0.3293 0.398 0.4093 ;
        RECT 0.398 0.0579 0.754 0.0973 ;
        RECT 0.754 0.0579 0.782 0.0973 ;
        RECT 0.754 0.0973 0.782 0.3293 ;
      LAYER V1 ;
        RECT 0.306 0.2253 0.334 0.244 ;
        RECT 0.306 0.4387 0.362 0.4573 ;
        RECT 0.498 0.2253 0.526 0.244 ;
      LAYER M1 ;
        RECT 0.08 0.108 0.099 0.1267 ;
        RECT 0.099 0.108 0.157 0.1267 ;
        RECT 0.099 0.328 0.157 0.3467 ;
        RECT 0.099 0.3467 0.157 0.384 ;
        RECT 0.157 0.108 0.306 0.1267 ;
        RECT 0.157 0.328 0.306 0.3467 ;
        RECT 0.306 0.108 0.334 0.1267 ;
        RECT 0.306 0.1267 0.334 0.328 ;
        RECT 0.306 0.328 0.334 0.3467 ;
        RECT 0.29 0.4387 0.434 0.4693 ;
        RECT 0.434 0.204 0.462 0.4387 ;
        RECT 0.434 0.4387 0.462 0.4693 ;
        RECT 0.498 0.1827 0.526 0.2853 ;
        RECT 0.37 0.0579 0.398 0.0973 ;
        RECT 0.37 0.0973 0.398 0.3293 ;
        RECT 0.37 0.3293 0.398 0.4093 ;
        RECT 0.398 0.0579 0.754 0.0973 ;
        RECT 0.754 0.0579 0.782 0.0973 ;
        RECT 0.754 0.0973 0.782 0.3293 ;
  END
END MUX2_X1_8T

MACRO NAND2_X1_8T
  CLASS core ;
  FOREIGN NAND2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3827 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3827 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0887 0.1419 0.128 ;
        RECT 0.114 0.128 0.1419 0.4253 ;
        RECT 0.1419 0.0887 0.176 0.128 ;
        RECT 0.176 0.0427 0.208 0.0887 ;
        RECT 0.176 0.0887 0.208 0.128 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END NAND2_X1_8T

MACRO NAND2_X2_8T
  CLASS core ;
  FOREIGN NAND2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.15 0.206 0.3687 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1827 0.078 0.4507 ;
        RECT 0.05 0.4507 0.078 0.4693 ;
        RECT 0.078 0.4507 0.306 0.4693 ;
        RECT 0.306 0.1827 0.334 0.4507 ;
        RECT 0.306 0.4507 0.334 0.4693 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.082 0.1419 0.1207 ;
        RECT 0.114 0.1207 0.1419 0.2827 ;
        RECT 0.114 0.2827 0.1419 0.398 ;
        RECT 0.114 0.398 0.1419 0.4267 ;
        RECT 0.1419 0.082 0.242 0.1207 ;
        RECT 0.1419 0.398 0.242 0.4267 ;
        RECT 0.242 0.082 0.27 0.1207 ;
        RECT 0.242 0.2827 0.27 0.398 ;
        RECT 0.242 0.398 0.27 0.4267 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NAND2_X2_8T

MACRO NAND3_X1_8T
  CLASS core ;
  FOREIGN NAND3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2133 0.27 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.17 0.206 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1433 0.078 0.3827 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.07334 0.0547 0.1419 0.0733 ;
        RECT 0.07334 0.0733 0.1419 0.1707 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
        RECT 0.114 0.3413 0.1419 0.4507 ;
        RECT 0.114 0.4507 0.1419 0.4693 ;
        RECT 0.1419 0.0547 0.242 0.0733 ;
        RECT 0.1419 0.4507 0.242 0.4693 ;
        RECT 0.242 0.0427 0.304 0.0547 ;
        RECT 0.242 0.0547 0.304 0.0733 ;
        RECT 0.242 0.4507 0.304 0.4693 ;
        RECT 0.304 0.0427 0.306 0.0547 ;
        RECT 0.304 0.0547 0.306 0.0733 ;
        RECT 0.304 0.0733 0.306 0.1707 ;
        RECT 0.304 0.4507 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.0547 ;
        RECT 0.306 0.0547 0.334 0.0733 ;
        RECT 0.306 0.0733 0.334 0.1707 ;
        RECT 0.306 0.3413 0.334 0.4507 ;
        RECT 0.306 0.4507 0.334 0.4693 ;
        RECT 0.334 0.0427 0.336 0.0547 ;
        RECT 0.334 0.0547 0.336 0.0733 ;
        RECT 0.334 0.0733 0.336 0.1707 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NAND3_X1_8T

MACRO NAND3_X2_8T
  CLASS core ;
  FOREIGN NAND3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.2133 0.526 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.301 0.166 0.339 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.027 0.3786 0.366 0.4173 ;
        RECT 0.366 0.3786 0.434 0.4173 ;
        RECT 0.434 0.124 0.462 0.3786 ;
        RECT 0.434 0.3786 0.462 0.4173 ;
        RECT 0.462 0.3786 0.494 0.4173 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.366 0.5307 ;
        RECT 0.366 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.074 0.498 0.0939 ;
        RECT 0.498 0.074 0.526 0.0939 ;
        RECT 0.498 0.0939 0.526 0.15 ;
        RECT 0.05 0.118 0.366 0.1393 ;
      LAYER M1 ;
        RECT 0.21 0.074 0.498 0.0939 ;
        RECT 0.498 0.074 0.526 0.0939 ;
        RECT 0.498 0.0939 0.526 0.15 ;
        RECT 0.05 0.118 0.366 0.1393 ;
  END
END NAND3_X2_8T

MACRO NAND4_X1_8T
  CLASS core ;
  FOREIGN NAND4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1707 0.398 0.3827 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.2987 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3827 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.3413 0.1419 0.43 ;
        RECT 0.114 0.43 0.1419 0.4693 ;
        RECT 0.1419 0.43 0.306 0.4693 ;
        RECT 0.306 0.1093 0.334 0.128 ;
        RECT 0.306 0.128 0.334 0.3413 ;
        RECT 0.306 0.3413 0.334 0.43 ;
        RECT 0.306 0.43 0.334 0.4693 ;
        RECT 0.334 0.1093 0.365 0.128 ;
        RECT 0.365 0.0427 0.403 0.1093 ;
        RECT 0.365 0.1093 0.403 0.128 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
END NAND4_X1_8T

MACRO NAND4_X2_8T
  CLASS core ;
  FOREIGN NAND4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.2387 0.594 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.2267 0.398 0.3507 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1613 0.206 0.3413 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1713 0.078 0.3413 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.37 0.144 0.384 ;
        RECT 0.112 0.384 0.144 0.4253 ;
        RECT 0.112 0.4253 0.144 0.444 ;
        RECT 0.144 0.4253 0.434 0.444 ;
        RECT 0.434 0.196 0.462 0.2147 ;
        RECT 0.434 0.2147 0.462 0.3653 ;
        RECT 0.434 0.3653 0.462 0.37 ;
        RECT 0.434 0.37 0.462 0.384 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.196 0.562 0.2147 ;
        RECT 0.462 0.3653 0.562 0.37 ;
        RECT 0.462 0.37 0.562 0.384 ;
        RECT 0.462 0.4253 0.562 0.444 ;
        RECT 0.562 0.196 0.59 0.2147 ;
        RECT 0.562 0.3653 0.59 0.37 ;
        RECT 0.562 0.37 0.59 0.384 ;
        RECT 0.562 0.384 0.59 0.4253 ;
        RECT 0.562 0.4253 0.59 0.444 ;
        RECT 0.59 0.196 0.654 0.2147 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.43 0.0867 ;
        RECT 0.274 0.1533 0.624 0.172 ;
        RECT 0.624 0.0427 0.656 0.1533 ;
        RECT 0.624 0.1533 0.656 0.172 ;
        RECT 0.146 0.1107 0.494 0.1293 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.43 0.0867 ;
        RECT 0.274 0.1533 0.624 0.172 ;
        RECT 0.624 0.0427 0.656 0.1533 ;
        RECT 0.624 0.1533 0.656 0.172 ;
        RECT 0.146 0.1107 0.494 0.1293 ;
  END
END NAND4_X2_8T

MACRO NOR2_X1_8T
  CLASS core ;
  FOREIGN NOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3413 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.384 ;
        RECT 0.114 0.384 0.1419 0.4233 ;
        RECT 0.1419 0.384 0.176 0.4233 ;
        RECT 0.176 0.384 0.208 0.4233 ;
        RECT 0.176 0.4233 0.208 0.4693 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.266 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.266 0.0187 ;
    END
  END VSS
END NOR2_X1_8T

MACRO NOR2_X2_8T
  CLASS core ;
  FOREIGN NOR2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1433 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.3293 ;
        RECT 0.078 0.0427 0.306 0.0613 ;
        RECT 0.306 0.0427 0.334 0.0613 ;
        RECT 0.306 0.0613 0.334 0.3293 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0853 0.1419 0.104 ;
        RECT 0.114 0.104 0.1419 0.2293 ;
        RECT 0.114 0.2293 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.0853 0.176 0.104 ;
        RECT 0.1419 0.3707 0.176 0.3893 ;
        RECT 0.176 0.0853 0.208 0.104 ;
        RECT 0.176 0.3707 0.208 0.3893 ;
        RECT 0.176 0.3893 0.208 0.4267 ;
        RECT 0.208 0.0853 0.242 0.104 ;
        RECT 0.242 0.0853 0.27 0.104 ;
        RECT 0.242 0.104 0.27 0.2293 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NOR2_X2_8T

MACRO NOR3_X1_8T
  CLASS core ;
  FOREIGN NOR3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2133 0.27 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1293 0.206 0.3687 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3687 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0427 0.1419 0.0613 ;
        RECT 0.114 0.0613 0.1419 0.1707 ;
        RECT 0.114 0.1707 0.1419 0.3413 ;
        RECT 0.114 0.3413 0.1419 0.4093 ;
        RECT 0.114 0.4093 0.1419 0.428 ;
        RECT 0.1419 0.0427 0.303 0.0613 ;
        RECT 0.1419 0.4093 0.303 0.428 ;
        RECT 0.303 0.0427 0.304 0.0613 ;
        RECT 0.303 0.0613 0.304 0.1707 ;
        RECT 0.303 0.4093 0.304 0.428 ;
        RECT 0.304 0.0427 0.336 0.0613 ;
        RECT 0.304 0.0613 0.336 0.1707 ;
        RECT 0.304 0.3413 0.336 0.4093 ;
        RECT 0.304 0.4093 0.336 0.428 ;
        RECT 0.304 0.428 0.336 0.4693 ;
        RECT 0.336 0.0427 0.337 0.0613 ;
        RECT 0.336 0.0613 0.337 0.1707 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
END NOR3_X1_8T

MACRO NOR3_X2_8T
  CLASS core ;
  FOREIGN NOR3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.1707 0.526 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.342 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.346 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0859 0.1027 0.434 0.1413 ;
        RECT 0.434 0.1027 0.462 0.1413 ;
        RECT 0.434 0.1413 0.462 0.384 ;
        RECT 0.462 0.1027 0.49 0.1413 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.526 0.5307 ;
        RECT 0.526 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.418 0.498 0.4367 ;
        RECT 0.498 0.344 0.526 0.418 ;
        RECT 0.498 0.418 0.526 0.4367 ;
        RECT 0.0859 0.3713 0.38 0.394 ;
      LAYER M1 ;
        RECT 0.21 0.418 0.498 0.4367 ;
        RECT 0.498 0.344 0.526 0.418 ;
        RECT 0.498 0.418 0.526 0.4367 ;
        RECT 0.0859 0.3713 0.38 0.394 ;
  END
END NOR3_X2_8T

MACRO NOR4_X1_8T
  CLASS core ;
  FOREIGN NOR4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1293 0.398 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1293 0.27 0.3413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.3827 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1293 0.078 0.3827 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.0427 0.1419 0.0679 ;
        RECT 0.114 0.0679 0.1419 0.1433 ;
        RECT 0.1419 0.0427 0.306 0.0679 ;
        RECT 0.306 0.0427 0.334 0.0679 ;
        RECT 0.306 0.0679 0.334 0.1433 ;
        RECT 0.306 0.1433 0.334 0.384 ;
        RECT 0.306 0.384 0.334 0.4027 ;
        RECT 0.334 0.384 0.365 0.4027 ;
        RECT 0.365 0.384 0.403 0.4027 ;
        RECT 0.365 0.4027 0.403 0.4693 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
END NOR4_X1_8T

MACRO NOR4_X2_8T
  CLASS core ;
  FOREIGN NOR4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.1707 0.594 0.2707 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.1613 0.398 0.292 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.3507 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.344 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.0679 0.144 0.0867 ;
        RECT 0.112 0.0867 0.144 0.128 ;
        RECT 0.112 0.128 0.144 0.142 ;
        RECT 0.144 0.0679 0.434 0.0867 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.128 0.462 0.142 ;
        RECT 0.434 0.142 0.462 0.1467 ;
        RECT 0.434 0.1467 0.462 0.2947 ;
        RECT 0.434 0.2947 0.462 0.3133 ;
        RECT 0.462 0.0679 0.562 0.0867 ;
        RECT 0.462 0.128 0.562 0.142 ;
        RECT 0.462 0.142 0.562 0.1467 ;
        RECT 0.462 0.2947 0.562 0.3133 ;
        RECT 0.562 0.0679 0.59 0.0867 ;
        RECT 0.562 0.0867 0.59 0.128 ;
        RECT 0.562 0.128 0.59 0.142 ;
        RECT 0.562 0.142 0.59 0.1467 ;
        RECT 0.562 0.2947 0.59 0.3133 ;
        RECT 0.59 0.2947 0.663 0.3133 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.43 0.5307 ;
        RECT 0.43 0.4933 0.494 0.5307 ;
        RECT 0.494 0.4933 0.656 0.5307 ;
        RECT 0.656 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.3799 0.494 0.4013 ;
        RECT 0.048 0.37 0.08 0.4253 ;
        RECT 0.048 0.4253 0.08 0.444 ;
        RECT 0.08 0.4253 0.43 0.444 ;
        RECT 0.338 0.3373 0.624 0.356 ;
        RECT 0.624 0.3373 0.656 0.356 ;
        RECT 0.624 0.356 0.656 0.4573 ;
      LAYER M1 ;
        RECT 0.21 0.3799 0.494 0.4013 ;
        RECT 0.048 0.37 0.08 0.4253 ;
        RECT 0.048 0.4253 0.08 0.444 ;
        RECT 0.08 0.4253 0.43 0.444 ;
        RECT 0.338 0.3373 0.624 0.356 ;
        RECT 0.624 0.3373 0.656 0.356 ;
        RECT 0.624 0.356 0.656 0.4573 ;
  END
END NOR4_X2_8T

MACRO OAI21_X1_8T
  CLASS core ;
  FOREIGN OAI21_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.1707 0.206 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.4227 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1707 0.334 0.384 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.424 ;
        RECT 0.114 0.424 0.1419 0.4453 ;
        RECT 0.1419 0.424 0.298 0.4453 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.0487 0.078 0.1033 ;
        RECT 0.05 0.1033 0.078 0.1247 ;
        RECT 0.078 0.1033 0.298 0.1247 ;
      LAYER M1 ;
        RECT 0.05 0.0487 0.078 0.1033 ;
        RECT 0.05 0.1033 0.078 0.1247 ;
        RECT 0.078 0.1033 0.298 0.1247 ;
  END
END OAI21_X1_8T

MACRO OAI21_X2_8T
  CLASS core ;
  FOREIGN OAI21_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.2133 0.403 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1613 0.1613 0.27 0.1886 ;
        RECT 0.242 0.1886 0.27 0.3347 ;
        RECT 0.242 0.3347 0.27 0.3533 ;
        RECT 0.27 0.3347 0.498 0.3533 ;
        RECT 0.498 0.1886 0.526 0.3347 ;
        RECT 0.498 0.3347 0.526 0.3533 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1707 0.1419 0.35 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.029 0.3799 0.178 0.4013 ;
        RECT 0.178 0.1107 0.206 0.1293 ;
        RECT 0.178 0.1293 0.206 0.1853 ;
        RECT 0.178 0.1853 0.206 0.3799 ;
        RECT 0.178 0.3799 0.206 0.4013 ;
        RECT 0.206 0.1107 0.426 0.1293 ;
        RECT 0.206 0.3799 0.426 0.4013 ;
        RECT 0.426 0.1107 0.434 0.1293 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.1853 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.498 0.0867 ;
        RECT 0.498 0.0679 0.526 0.0867 ;
        RECT 0.498 0.0867 0.526 0.142 ;
        RECT 0.498 0.142 0.526 0.1433 ;
        RECT 0.146 0.4253 0.535 0.444 ;
      LAYER M1 ;
        RECT 0.048 0.0679 0.08 0.0867 ;
        RECT 0.048 0.0867 0.08 0.142 ;
        RECT 0.08 0.0679 0.498 0.0867 ;
        RECT 0.498 0.0679 0.526 0.0867 ;
        RECT 0.498 0.0867 0.526 0.142 ;
        RECT 0.498 0.142 0.526 0.1433 ;
        RECT 0.146 0.4253 0.535 0.444 ;
  END
END OAI21_X2_8T

MACRO OAI22_X1_8T
  CLASS core ;
  FOREIGN OAI22_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.1327 0.27 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.186 0.398 0.384 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.128 0.206 0.3413 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.128 0.08 0.384 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.4253 0.306 0.444 ;
        RECT 0.306 0.1213 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.444 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.0673 0.37 0.0873 ;
        RECT 0.37 0.0673 0.398 0.0873 ;
        RECT 0.37 0.0873 0.398 0.1407 ;
      LAYER M1 ;
        RECT 0.05 0.0673 0.37 0.0873 ;
        RECT 0.37 0.0673 0.398 0.0873 ;
        RECT 0.37 0.0873 0.398 0.1407 ;
  END
END OAI22_X1_8T

MACRO OAI22_X2_8T
  CLASS core ;
  FOREIGN OAI22_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.1707 0.462 0.186 ;
        RECT 0.434 0.186 0.462 0.3107 ;
        RECT 0.434 0.3107 0.462 0.3293 ;
        RECT 0.462 0.3107 0.6899 0.3293 ;
        RECT 0.6899 0.186 0.718 0.3107 ;
        RECT 0.6899 0.3107 0.718 0.3293 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.1707 0.59 0.2653 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.1613 0.334 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3413 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2573 0.27 0.3533 ;
        RECT 0.242 0.3533 0.27 0.372 ;
        RECT 0.27 0.3533 0.37 0.372 ;
        RECT 0.37 0.1127 0.398 0.1313 ;
        RECT 0.37 0.1313 0.398 0.1853 ;
        RECT 0.37 0.1853 0.398 0.2573 ;
        RECT 0.37 0.2573 0.398 0.3533 ;
        RECT 0.37 0.3533 0.398 0.372 ;
        RECT 0.398 0.1127 0.626 0.1313 ;
        RECT 0.398 0.3533 0.626 0.372 ;
        RECT 0.626 0.1127 0.654 0.1313 ;
        RECT 0.626 0.1313 0.654 0.1853 ;
        RECT 0.626 0.3533 0.654 0.372 ;
        RECT 0.654 0.3533 0.6899 0.372 ;
        RECT 0.6899 0.3533 0.718 0.372 ;
        RECT 0.6899 0.372 0.718 0.448 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.362 0.5307 ;
        RECT 0.362 0.4933 0.654 0.5307 ;
        RECT 0.654 0.4933 0.718 0.5307 ;
        RECT 0.718 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.402 0.4027 0.626 0.424 ;
        RECT 0.626 0.4027 0.654 0.424 ;
        RECT 0.626 0.424 0.654 0.4639 ;
        RECT 0.041 0.066 0.6899 0.0887 ;
        RECT 0.6899 0.066 0.718 0.0887 ;
        RECT 0.6899 0.0887 0.718 0.1407 ;
        RECT 0.05 0.408 0.362 0.4467 ;
      LAYER M1 ;
        RECT 0.402 0.4027 0.626 0.424 ;
        RECT 0.626 0.4027 0.654 0.424 ;
        RECT 0.626 0.424 0.654 0.4639 ;
        RECT 0.041 0.066 0.6899 0.0887 ;
        RECT 0.6899 0.066 0.718 0.0887 ;
        RECT 0.6899 0.0887 0.718 0.1407 ;
        RECT 0.05 0.408 0.362 0.4467 ;
  END
END OAI22_X2_8T

MACRO OR2_X1_8T
  CLASS core ;
  FOREIGN OR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.064 0.206 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.162 0.078 0.4273 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.076 0.334 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.394 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.394 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.224 ;
        RECT 0.114 0.224 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.3707 0.242 0.3893 ;
        RECT 0.242 0.224 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
      LAYER M1 ;
        RECT 0.114 0.0867 0.1419 0.224 ;
        RECT 0.114 0.224 0.1419 0.3707 ;
        RECT 0.114 0.3707 0.1419 0.3893 ;
        RECT 0.1419 0.3707 0.242 0.3893 ;
        RECT 0.242 0.224 0.27 0.3707 ;
        RECT 0.242 0.3707 0.27 0.3893 ;
  END
END OR2_X1_8T

MACRO OR2_X2_8T
  CLASS core ;
  FOREIGN OR2_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1613 0.1419 0.3413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3413 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.0427 0.306 0.09 ;
        RECT 0.302 0.4253 0.306 0.4693 ;
        RECT 0.306 0.0427 0.334 0.09 ;
        RECT 0.306 0.09 0.334 0.4253 ;
        RECT 0.306 0.4253 0.334 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.27 0.5307 ;
        RECT 0.27 0.4933 0.458 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.458 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.077 0.1027 0.146 0.1253 ;
        RECT 0.146 0.1027 0.242 0.1253 ;
        RECT 0.146 0.3867 0.242 0.4053 ;
        RECT 0.242 0.1027 0.27 0.1253 ;
        RECT 0.242 0.1253 0.27 0.3867 ;
        RECT 0.242 0.3867 0.27 0.4053 ;
      LAYER M1 ;
        RECT 0.077 0.1027 0.146 0.1253 ;
        RECT 0.146 0.1027 0.242 0.1253 ;
        RECT 0.146 0.3867 0.242 0.4053 ;
        RECT 0.242 0.1027 0.27 0.1253 ;
        RECT 0.242 0.1253 0.27 0.3867 ;
        RECT 0.242 0.3867 0.27 0.4053 ;
  END
END OR2_X2_8T

MACRO OR3_X1_8T
  CLASS core ;
  FOREIGN OR3_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.128 0.208 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.128 0.083 0.384 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.076 0.462 0.436 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.234 0.5307 ;
        RECT 0.234 0.4933 0.398 0.5307 ;
        RECT 0.398 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.0727 0.278 0.0913 ;
        RECT 0.278 0.0727 0.37 0.0913 ;
        RECT 0.278 0.4207 0.37 0.4487 ;
        RECT 0.37 0.0727 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4487 ;
        RECT 0.0859 0.424 0.234 0.4453 ;
      LAYER M1 ;
        RECT 0.054 0.0727 0.278 0.0913 ;
        RECT 0.278 0.0727 0.37 0.0913 ;
        RECT 0.278 0.4207 0.37 0.4487 ;
        RECT 0.37 0.0727 0.398 0.0913 ;
        RECT 0.37 0.0913 0.398 0.4207 ;
        RECT 0.37 0.4207 0.398 0.4487 ;
        RECT 0.0859 0.424 0.234 0.4453 ;
  END
END OR3_X1_8T

MACRO OR3_X2_8T
  CLASS core ;
  FOREIGN OR3_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.17 0.1419 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1707 0.078 0.3507 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.154 0.27 0.2987 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.0427 0.37 0.0867 ;
        RECT 0.366 0.424 0.37 0.4693 ;
        RECT 0.37 0.0427 0.398 0.0867 ;
        RECT 0.37 0.0867 0.398 0.424 ;
        RECT 0.37 0.424 0.398 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.302 0.5307 ;
        RECT 0.302 0.4933 0.334 0.5307 ;
        RECT 0.334 0.4933 0.522 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.522 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.3819 0.078 0.402 ;
        RECT 0.05 0.402 0.078 0.4573 ;
        RECT 0.078 0.3819 0.302 0.402 ;
        RECT 0.06 0.1033 0.1409 0.1247 ;
        RECT 0.1409 0.1033 0.306 0.1247 ;
        RECT 0.1409 0.3367 0.306 0.358 ;
        RECT 0.306 0.1033 0.334 0.1247 ;
        RECT 0.306 0.1247 0.334 0.3367 ;
        RECT 0.306 0.3367 0.334 0.358 ;
      LAYER M1 ;
        RECT 0.05 0.3819 0.078 0.402 ;
        RECT 0.05 0.402 0.078 0.4573 ;
        RECT 0.078 0.3819 0.302 0.402 ;
        RECT 0.06 0.1033 0.1409 0.1247 ;
        RECT 0.1409 0.1033 0.306 0.1247 ;
        RECT 0.1409 0.3367 0.306 0.358 ;
        RECT 0.306 0.1033 0.334 0.1247 ;
        RECT 0.306 0.1247 0.334 0.3367 ;
        RECT 0.306 0.3367 0.334 0.358 ;
  END
END OR3_X2_8T

MACRO OR4_X1_8T
  CLASS core ;
  FOREIGN OR4_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.128 0.398 0.384 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.128 0.272 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.132 0.1419 0.384 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.128 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.076 0.526 0.4267 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.298 0.5307 ;
        RECT 0.298 0.4933 0.462 0.5307 ;
        RECT 0.462 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.0679 0.338 0.0867 ;
        RECT 0.338 0.0679 0.434 0.0867 ;
        RECT 0.338 0.42 0.434 0.4413 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.42 ;
        RECT 0.434 0.42 0.462 0.4413 ;
        RECT 0.146 0.4113 0.298 0.4367 ;
      LAYER M1 ;
        RECT 0.054 0.0679 0.338 0.0867 ;
        RECT 0.338 0.0679 0.434 0.0867 ;
        RECT 0.338 0.42 0.434 0.4413 ;
        RECT 0.434 0.0679 0.462 0.0867 ;
        RECT 0.434 0.0867 0.462 0.42 ;
        RECT 0.434 0.42 0.462 0.4413 ;
        RECT 0.146 0.4113 0.298 0.4367 ;
  END
END OR4_X1_8T

MACRO OR4_X2_8T
  CLASS core ;
  FOREIGN OR4_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.128 0.334 0.3533 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.142 0.27 0.384 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.142 0.1419 0.384 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1273 0.078 0.384 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.0853 0.528 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.302 0.5307 ;
        RECT 0.302 0.4933 0.46 0.5307 ;
        RECT 0.46 0.4933 0.65 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.65 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.4153 0.302 0.454 ;
        RECT 0.054 0.0579 0.342 0.0967 ;
        RECT 0.342 0.0579 0.432 0.0967 ;
        RECT 0.342 0.3786 0.432 0.416 ;
        RECT 0.432 0.0579 0.46 0.0967 ;
        RECT 0.432 0.0967 0.46 0.3786 ;
        RECT 0.432 0.3786 0.46 0.416 ;
      LAYER M1 ;
        RECT 0.146 0.4153 0.302 0.454 ;
        RECT 0.054 0.0579 0.342 0.0967 ;
        RECT 0.342 0.0579 0.432 0.0967 ;
        RECT 0.342 0.3786 0.432 0.416 ;
        RECT 0.432 0.0579 0.46 0.0967 ;
        RECT 0.432 0.0967 0.46 0.3786 ;
        RECT 0.432 0.3786 0.46 0.416 ;
  END
END OR4_X2_8T

MACRO SDFFRNQ_X1_8T
  CLASS core ;
  FOREIGN SDFFRNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.242 0.515 0.352 ;
        RECT 0.515 0.242 0.526 0.352 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.965 0.2253 1.454 0.244 ;
        RECT 1.454 0.2253 1.592 0.244 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.248 0.334 0.3813 ;
        RECT 0.306 0.3813 0.334 0.4 ;
        RECT 0.334 0.3813 0.515 0.4 ;
        RECT 0.515 0.3813 0.562 0.4 ;
        RECT 0.562 0.2093 0.59 0.248 ;
        RECT 0.562 0.248 0.59 0.3813 ;
        RECT 0.562 0.3813 0.59 0.4 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.3413 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.184 0.078 0.356 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.0427 1.872 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.754 0.5307 ;
        RECT 0.754 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 1.066 0.5307 ;
        RECT 1.066 0.4933 1.422 0.5307 ;
        RECT 1.422 0.4933 1.49 0.5307 ;
        RECT 1.49 0.4933 1.742 0.5307 ;
        RECT 1.742 0.4933 1.93 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.93 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.121 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.121 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER M1 ;
        RECT 0.045 0.064 0.083 0.1359 ;
        RECT 0.045 0.1359 0.083 0.1547 ;
        RECT 0.045 0.4027 0.083 0.4213 ;
        RECT 0.045 0.4213 0.083 0.4586 ;
        RECT 0.083 0.1359 0.114 0.1547 ;
        RECT 0.083 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1359 0.1419 0.1547 ;
        RECT 0.114 0.1547 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.064 0.27 0.178 ;
        RECT 0.242 0.178 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.448 ;
        RECT 0.27 0.178 0.515 0.1967 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.754 0.4453 ;
        RECT 0.754 0.1647 0.782 0.364 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 1.061 0.16 1.098 0.2973 ;
        RECT 1.202 0.114 1.23 0.3407 ;
        RECT 1.458 0.0973 1.49 0.4653 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0427 1.358 0.0613 ;
        RECT 1.33 0.0613 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0427 1.607 0.0613 ;
        RECT 1.607 0.0427 1.635 0.0613 ;
        RECT 1.607 0.0613 1.635 0.244 ;
        RECT 1.554 0.3067 1.582 0.416 ;
        RECT 1.554 0.416 1.582 0.4533 ;
        RECT 1.582 0.416 1.714 0.4533 ;
        RECT 1.714 0.048 1.742 0.3067 ;
        RECT 1.714 0.3067 1.742 0.416 ;
        RECT 1.714 0.416 1.742 0.4533 ;
        RECT 0.178 0.0833 0.206 0.3827 ;
        RECT 0.6899 0.258 0.718 0.3933 ;
        RECT 0.8179 0.1713 0.85 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 0.991 0.1613 1.025 0.2813 ;
        RECT 0.79 0.424 1.066 0.4453 ;
        RECT 0.904 0.1827 0.932 0.3267 ;
        RECT 0.904 0.3267 0.932 0.3453 ;
        RECT 0.932 0.3267 1.1339 0.3453 ;
        RECT 1.1339 0.0547 1.166 0.1827 ;
        RECT 1.1339 0.1827 1.166 0.3267 ;
        RECT 1.1339 0.3267 1.166 0.3453 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.3293 ;
        RECT 1.532 0.1027 1.571 0.2773 ;
      LAYER V1 ;
        RECT 0.114 0.1827 0.1419 0.2013 ;
        RECT 0.178 0.3533 0.206 0.372 ;
        RECT 0.6899 0.3533 0.718 0.372 ;
        RECT 0.754 0.268 0.782 0.2867 ;
        RECT 0.8179 0.1827 0.846 0.2013 ;
        RECT 0.997 0.2253 1.025 0.244 ;
        RECT 1.061 0.268 1.089 0.2867 ;
        RECT 1.202 0.1827 1.23 0.2013 ;
        RECT 1.266 0.3533 1.294 0.372 ;
        RECT 1.3939 0.1827 1.422 0.2013 ;
        RECT 1.532 0.2253 1.56 0.244 ;
      LAYER M1 ;
        RECT 0.045 0.064 0.083 0.1359 ;
        RECT 0.045 0.1359 0.083 0.1547 ;
        RECT 0.045 0.4027 0.083 0.4213 ;
        RECT 0.045 0.4213 0.083 0.4586 ;
        RECT 0.083 0.1359 0.114 0.1547 ;
        RECT 0.083 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1359 0.1419 0.1547 ;
        RECT 0.114 0.1547 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.064 0.27 0.178 ;
        RECT 0.242 0.178 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.448 ;
        RECT 0.27 0.178 0.515 0.1967 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.754 0.4453 ;
        RECT 0.754 0.1647 0.782 0.364 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 1.061 0.16 1.098 0.2973 ;
        RECT 1.202 0.114 1.23 0.3407 ;
        RECT 1.458 0.0973 1.49 0.4653 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0427 1.358 0.0613 ;
        RECT 1.33 0.0613 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0427 1.607 0.0613 ;
        RECT 1.607 0.0427 1.635 0.0613 ;
        RECT 1.607 0.0613 1.635 0.244 ;
        RECT 1.554 0.3067 1.582 0.416 ;
        RECT 1.554 0.416 1.582 0.4533 ;
        RECT 1.582 0.416 1.714 0.4533 ;
        RECT 1.714 0.048 1.742 0.3067 ;
        RECT 1.714 0.3067 1.742 0.416 ;
        RECT 1.714 0.416 1.742 0.4533 ;
        RECT 0.178 0.0833 0.206 0.3827 ;
        RECT 0.6899 0.258 0.718 0.3933 ;
        RECT 0.8179 0.1713 0.85 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 0.991 0.1613 1.025 0.2813 ;
        RECT 0.79 0.424 1.066 0.4453 ;
        RECT 0.904 0.1827 0.932 0.3267 ;
        RECT 0.904 0.3267 0.932 0.3453 ;
        RECT 0.932 0.3267 1.1339 0.3453 ;
        RECT 1.1339 0.0547 1.166 0.1827 ;
        RECT 1.1339 0.1827 1.166 0.3267 ;
        RECT 1.1339 0.3267 1.166 0.3453 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.3293 ;
        RECT 1.532 0.1027 1.571 0.2773 ;
  END
END SDFFRNQ_X1_8T

MACRO SDFFSNQ_X1_8T
  CLASS core ;
  FOREIGN SDFFSNQ_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.512 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.256 0.51 0.352 ;
        RECT 0.51 0.256 0.526 0.352 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.248 0.334 0.3813 ;
        RECT 0.306 0.3813 0.334 0.4 ;
        RECT 0.334 0.3813 0.51 0.4 ;
        RECT 0.51 0.3813 0.562 0.4 ;
        RECT 0.562 0.2093 0.59 0.248 ;
        RECT 0.562 0.248 0.59 0.3813 ;
        RECT 0.562 0.3813 0.59 0.4 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.3413 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.958 0.2253 1.454 0.244 ;
        RECT 1.454 0.2253 1.586 0.244 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1813 0.078 0.3413 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.0427 1.872 0.4693 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.206 0.5307 ;
        RECT 0.206 0.4933 0.49336 0.5307 ;
        RECT 0.49336 0.4933 0.782 0.5307 ;
        RECT 0.782 0.4933 0.862 0.5307 ;
        RECT 0.862 0.4933 1.646 0.5307 ;
        RECT 1.646 0.4933 1.742 0.5307 ;
        RECT 1.742 0.4933 1.93 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.93 0.0187 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.114 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER MINT1 ;
        RECT 0.146 0.3533 1.326 0.372 ;
        RECT 0.722 0.268 1.114 0.2867 ;
        RECT 0.082 0.1827 1.454 0.2013 ;
      LAYER M1 ;
        RECT 0.048 0.0427 0.08 0.1333 ;
        RECT 0.048 0.1333 0.08 0.133328 ;
        RECT 0.048 0.4027 0.08 0.4213 ;
        RECT 0.048 0.4213 0.08 0.4586 ;
        RECT 0.08 0.1333 0.114 0.133328 ;
        RECT 0.08 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1333 0.1419 0.133328 ;
        RECT 0.114 0.152 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.0547 0.27 0.1773 ;
        RECT 0.242 0.1773 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.1973 ;
        RECT 0.242 0.1973 0.27 0.4573 ;
        RECT 0.27 0.1773 0.434 0.1967 ;
        RECT 0.434 0.1773 0.51 0.1967 ;
        RECT 0.434 0.1967 0.51 0.1973 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.746 0.4453 ;
        RECT 0.754 0.1587 0.782 0.3647 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 0.98 0.2147 1.018 0.2793 ;
        RECT 0.898 0.1827 0.926 0.3247 ;
        RECT 0.898 0.3247 0.926 0.3433 ;
        RECT 0.926 0.3247 1.008 0.3433 ;
        RECT 1.008 0.3247 1.04 0.3433 ;
        RECT 1.008 0.3433 1.04 0.4693 ;
        RECT 1.04 0.3247 1.1379 0.3433 ;
        RECT 1.1379 0.0653 1.166 0.1827 ;
        RECT 1.1379 0.1827 1.166 0.3247 ;
        RECT 1.1379 0.3247 1.166 0.3433 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.268 ;
        RECT 1.526 0.1227 1.554 0.2687 ;
        RECT 1.402 0.4253 1.646 0.444 ;
        RECT 0.178 0.064 0.206 0.4127 ;
        RECT 0.654 0.258 0.682 0.3827 ;
        RECT 0.83 0.1713 0.862 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 1.054 0.16 1.092 0.2973 ;
        RECT 1.202 0.114 1.23 0.2553 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0547 1.358 0.0733 ;
        RECT 1.33 0.0733 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0547 1.607 0.0733 ;
        RECT 1.607 0.0547 1.645 0.0733 ;
        RECT 1.607 0.0733 1.645 0.244 ;
        RECT 1.462 0.268 1.49 0.3827 ;
        RECT 1.462 0.3827 1.49 0.4013 ;
        RECT 1.49 0.3827 1.714 0.4013 ;
        RECT 1.714 0.064 1.742 0.268 ;
        RECT 1.714 0.268 1.742 0.3827 ;
        RECT 1.714 0.3827 1.742 0.4013 ;
      LAYER V1 ;
        RECT 0.114 0.1827 0.1419 0.2013 ;
        RECT 0.178 0.3533 0.206 0.372 ;
        RECT 0.654 0.3533 0.682 0.372 ;
        RECT 0.754 0.268 0.782 0.2867 ;
        RECT 0.834 0.1827 0.862 0.2013 ;
        RECT 0.99 0.2253 1.018 0.244 ;
        RECT 1.054 0.268 1.082 0.2867 ;
        RECT 1.202 0.1827 1.23 0.2013 ;
        RECT 1.266 0.3533 1.294 0.372 ;
        RECT 1.3939 0.1827 1.422 0.2013 ;
        RECT 1.526 0.2253 1.554 0.244 ;
      LAYER M1 ;
        RECT 0.048 0.0427 0.08 0.1333 ;
        RECT 0.048 0.1333 0.08 0.133328 ;
        RECT 0.048 0.4027 0.08 0.4213 ;
        RECT 0.048 0.4213 0.08 0.4586 ;
        RECT 0.08 0.1333 0.114 0.133328 ;
        RECT 0.08 0.4027 0.114 0.4213 ;
        RECT 0.114 0.1333 0.1419 0.133328 ;
        RECT 0.114 0.152 0.1419 0.4027 ;
        RECT 0.114 0.4027 0.1419 0.4213 ;
        RECT 0.242 0.0547 0.27 0.1773 ;
        RECT 0.242 0.1773 0.27 0.1967 ;
        RECT 0.242 0.1967 0.27 0.1973 ;
        RECT 0.242 0.1973 0.27 0.4573 ;
        RECT 0.27 0.1773 0.434 0.1967 ;
        RECT 0.434 0.1773 0.51 0.1967 ;
        RECT 0.434 0.1967 0.51 0.1973 ;
        RECT 0.338 0.1227 0.626 0.1413 ;
        RECT 0.626 0.1227 0.654 0.1413 ;
        RECT 0.626 0.1413 0.654 0.184 ;
        RECT 0.392 0.424 0.746 0.4453 ;
        RECT 0.754 0.1587 0.782 0.3647 ;
        RECT 0.466 0.0679 0.878 0.0867 ;
        RECT 0.98 0.2147 1.018 0.2793 ;
        RECT 0.898 0.1827 0.926 0.3247 ;
        RECT 0.898 0.3247 0.926 0.3433 ;
        RECT 0.926 0.3247 1.008 0.3433 ;
        RECT 1.008 0.3247 1.04 0.3433 ;
        RECT 1.008 0.3433 1.04 0.4693 ;
        RECT 1.04 0.3247 1.1379 0.3433 ;
        RECT 1.1379 0.0653 1.166 0.1827 ;
        RECT 1.1379 0.1827 1.166 0.3247 ;
        RECT 1.1379 0.3247 1.166 0.3433 ;
        RECT 1.266 0.1187 1.294 0.3827 ;
        RECT 1.3939 0.1187 1.422 0.268 ;
        RECT 1.526 0.1227 1.554 0.2687 ;
        RECT 1.402 0.4253 1.646 0.444 ;
        RECT 0.178 0.064 0.206 0.4127 ;
        RECT 0.654 0.258 0.682 0.3827 ;
        RECT 0.83 0.1713 0.862 0.3127 ;
        RECT 0.6899 0.1107 0.718 0.1293 ;
        RECT 0.6899 0.1293 0.718 0.184 ;
        RECT 0.718 0.1107 0.942 0.1293 ;
        RECT 1.054 0.16 1.092 0.2973 ;
        RECT 1.202 0.114 1.23 0.2553 ;
        RECT 1.165 0.412 1.33 0.4307 ;
        RECT 1.33 0.0547 1.358 0.0733 ;
        RECT 1.33 0.0733 1.358 0.244 ;
        RECT 1.33 0.244 1.358 0.412 ;
        RECT 1.33 0.412 1.358 0.4307 ;
        RECT 1.358 0.0547 1.607 0.0733 ;
        RECT 1.607 0.0547 1.645 0.0733 ;
        RECT 1.607 0.0733 1.645 0.244 ;
        RECT 1.462 0.268 1.49 0.3827 ;
        RECT 1.462 0.3827 1.49 0.4013 ;
        RECT 1.49 0.3827 1.714 0.4013 ;
        RECT 1.714 0.064 1.742 0.268 ;
        RECT 1.714 0.268 1.742 0.3827 ;
        RECT 1.714 0.3827 1.742 0.4013 ;
  END
END SDFFSNQ_X1_8T

MACRO TBUF_X1_8T
  CLASS core ;
  FOREIGN TBUF_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.3467 ;
        RECT 0.1419 0.328 0.206 0.3467 ;
        RECT 0.206 0.328 0.242 0.3467 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.328 ;
        RECT 0.242 0.328 0.27 0.3467 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2467 0.462 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.0427 0.656 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.588 0.5307 ;
        RECT 0.588 0.4933 0.714 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.714 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2787 ;
        RECT 0.05 0.2787 0.078 0.4573 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2787 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.51 0.0867 ;
        RECT 0.51 0.0679 0.542 0.0867 ;
        RECT 0.51 0.0867 0.542 0.1533 ;
        RECT 0.51 0.1533 0.542 0.172 ;
        RECT 0.51 0.172 0.542 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2507 ;
        RECT 0.37 0.2507 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.56 0.444 ;
        RECT 0.56 0.2507 0.588 0.4253 ;
        RECT 0.56 0.4253 0.588 0.444 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2787 ;
        RECT 0.05 0.2787 0.078 0.4573 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2787 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.51 0.0867 ;
        RECT 0.51 0.0679 0.542 0.0867 ;
        RECT 0.51 0.0867 0.542 0.1533 ;
        RECT 0.51 0.1533 0.542 0.172 ;
        RECT 0.51 0.172 0.542 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2507 ;
        RECT 0.37 0.2507 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.56 0.444 ;
        RECT 0.56 0.2507 0.588 0.4253 ;
        RECT 0.56 0.4253 0.588 0.444 ;
  END
END TBUF_X1_8T

MACRO TBUF_X2_8T
  CLASS core ;
  FOREIGN TBUF_X2_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.3547 ;
        RECT 0.1419 0.336 0.206 0.3547 ;
        RECT 0.206 0.336 0.242 0.3547 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.336 ;
        RECT 0.242 0.336 0.27 0.3547 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2547 0.462 0.384 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.0467 0.656 0.4639 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.53 0.5307 ;
        RECT 0.53 0.4933 0.778 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.778 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.408 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.482 0.0867 ;
        RECT 0.482 0.0679 0.514 0.0867 ;
        RECT 0.482 0.0867 0.514 0.1533 ;
        RECT 0.482 0.1533 0.514 0.172 ;
        RECT 0.482 0.172 0.514 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2953 ;
        RECT 0.37 0.2953 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.498 0.444 ;
        RECT 0.498 0.2953 0.53 0.4253 ;
        RECT 0.498 0.4253 0.53 0.444 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.408 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.2093 ;
        RECT 0.306 0.2093 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.482 0.0867 ;
        RECT 0.482 0.0679 0.514 0.0867 ;
        RECT 0.482 0.0867 0.514 0.1533 ;
        RECT 0.482 0.1533 0.514 0.172 ;
        RECT 0.482 0.172 0.514 0.2093 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2953 ;
        RECT 0.37 0.2953 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.498 0.444 ;
        RECT 0.498 0.2953 0.53 0.4253 ;
        RECT 0.498 0.4253 0.53 0.444 ;
  END
END TBUF_X2_8T

MACRO TBUF_X4_8T
  CLASS core ;
  FOREIGN TBUF_X4_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.3227 ;
        RECT 0.114 0.3227 0.1419 0.3413 ;
        RECT 0.1419 0.3227 0.206 0.3413 ;
        RECT 0.206 0.3227 0.242 0.3413 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.3227 ;
        RECT 0.242 0.3227 0.27 0.3413 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.2306 0.462 0.396 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6879 0.0427 0.72 0.1493 ;
        RECT 0.6879 0.1493 0.72 0.1707 ;
        RECT 0.6879 0.3413 0.72 0.36 ;
        RECT 0.6879 0.36 0.72 0.3806 ;
        RECT 0.6879 0.3806 0.72 0.4693 ;
        RECT 0.72 0.1493 0.8129 0.1707 ;
        RECT 0.72 0.3413 0.8129 0.36 ;
        RECT 0.8129 0.0427 0.8139 0.1493 ;
        RECT 0.8129 0.1493 0.8139 0.1707 ;
        RECT 0.8129 0.3413 0.8139 0.36 ;
        RECT 0.8139 0.0427 0.8159 0.1493 ;
        RECT 0.8139 0.1493 0.8159 0.1707 ;
        RECT 0.8139 0.3413 0.8159 0.36 ;
        RECT 0.8159 0.0427 0.838 0.1493 ;
        RECT 0.8159 0.1493 0.838 0.1707 ;
        RECT 0.8159 0.3413 0.838 0.36 ;
        RECT 0.8159 0.36 0.838 0.3806 ;
        RECT 0.8159 0.3806 0.838 0.4693 ;
        RECT 0.838 0.0427 0.848 0.1493 ;
        RECT 0.838 0.1493 0.848 0.1707 ;
        RECT 0.838 0.3413 0.848 0.36 ;
        RECT 0.838 0.36 0.848 0.3806 ;
        RECT 0.838 0.3806 0.848 0.4693 ;
        RECT 0.848 0.0427 0.851 0.1493 ;
        RECT 0.848 0.1493 0.851 0.1707 ;
        RECT 0.848 0.3413 0.851 0.36 ;
        RECT 0.848 0.36 0.851 0.3806 ;
        RECT 0.851 0.1493 0.882 0.1707 ;
        RECT 0.851 0.3413 0.882 0.36 ;
        RECT 0.851 0.36 0.882 0.3806 ;
        RECT 0.882 0.1493 0.91 0.1707 ;
        RECT 0.882 0.1707 0.91 0.3413 ;
        RECT 0.882 0.3413 0.91 0.36 ;
        RECT 0.882 0.36 0.91 0.3806 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.8139 0.5307 ;
        RECT 0.8139 0.4933 0.838 0.5307 ;
        RECT 0.838 0.4933 0.97 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.97 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2587 ;
        RECT 0.37 0.2587 0.398 0.276 ;
        RECT 0.37 0.276 0.398 0.3053 ;
        RECT 0.37 0.3053 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.526 0.444 ;
        RECT 0.526 0.2587 0.582 0.276 ;
        RECT 0.526 0.276 0.582 0.3053 ;
        RECT 0.526 0.3053 0.582 0.4253 ;
        RECT 0.526 0.4253 0.582 0.444 ;
        RECT 0.582 0.276 0.8139 0.3053 ;
        RECT 0.05 0.064 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.396 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.1947 ;
        RECT 0.306 0.1947 0.334 0.2133 ;
        RECT 0.306 0.2133 0.334 0.2347 ;
        RECT 0.306 0.2347 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.526 0.0867 ;
        RECT 0.526 0.0679 0.582 0.0867 ;
        RECT 0.526 0.0867 0.582 0.1533 ;
        RECT 0.526 0.1533 0.582 0.172 ;
        RECT 0.526 0.172 0.582 0.1947 ;
        RECT 0.526 0.1947 0.582 0.2133 ;
        RECT 0.526 0.2133 0.582 0.2347 ;
        RECT 0.582 0.1947 0.838 0.2133 ;
      LAYER M1 ;
        RECT 0.082 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2587 ;
        RECT 0.37 0.2587 0.398 0.276 ;
        RECT 0.37 0.276 0.398 0.3053 ;
        RECT 0.37 0.3053 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.526 0.444 ;
        RECT 0.526 0.2587 0.582 0.276 ;
        RECT 0.526 0.276 0.582 0.3053 ;
        RECT 0.526 0.3053 0.582 0.4253 ;
        RECT 0.526 0.4253 0.582 0.444 ;
        RECT 0.582 0.276 0.8139 0.3053 ;
        RECT 0.05 0.064 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.396 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.146 0.3786 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3786 0.23 0.4013 ;
        RECT 0.23 0.0679 0.306 0.0867 ;
        RECT 0.1533 0.1533 0.306 0.172 ;
        RECT 0.23 0.3786 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.172 ;
        RECT 0.306 0.172 0.334 0.1947 ;
        RECT 0.306 0.1947 0.334 0.2133 ;
        RECT 0.306 0.2133 0.334 0.2347 ;
        RECT 0.306 0.2347 0.334 0.3786 ;
        RECT 0.306 0.3786 0.334 0.4013 ;
        RECT 0.334 0.0679 0.526 0.0867 ;
        RECT 0.526 0.0679 0.582 0.0867 ;
        RECT 0.526 0.0867 0.582 0.1533 ;
        RECT 0.526 0.1533 0.582 0.172 ;
        RECT 0.526 0.172 0.582 0.1947 ;
        RECT 0.526 0.1947 0.582 0.2133 ;
        RECT 0.526 0.2133 0.582 0.2347 ;
        RECT 0.582 0.1947 0.838 0.2133 ;
  END
END TBUF_X4_8T

MACRO TBUF_X8_8T
  CLASS core ;
  FOREIGN TBUF_X8_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.3227 ;
        RECT 0.114 0.3227 0.1419 0.3413 ;
        RECT 0.1419 0.3227 0.222 0.3413 ;
        RECT 0.222 0.3227 0.306 0.3413 ;
        RECT 0.306 0.2133 0.334 0.256 ;
        RECT 0.306 0.256 0.334 0.3227 ;
        RECT 0.306 0.3227 0.334 0.3413 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.2306 0.526 0.268 ;
        RECT 0.498 0.268 0.526 0.2893 ;
        RECT 0.498 0.2893 0.526 0.384 ;
        RECT 0.526 0.268 0.622 0.2893 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8159 0.0427 0.848 0.0887 ;
        RECT 0.8159 0.0887 0.848 0.1067 ;
        RECT 0.8159 0.1067 0.848 0.128 ;
        RECT 0.8159 0.346 0.848 0.3847 ;
        RECT 0.8159 0.3847 0.848 0.3853 ;
        RECT 0.8159 0.3853 0.848 0.4693 ;
        RECT 0.848 0.1067 1.183 0.128 ;
        RECT 0.848 0.346 1.183 0.3847 ;
        RECT 1.183 0.1067 1.198 0.128 ;
        RECT 1.183 0.346 1.198 0.3847 ;
        RECT 1.198 0.1067 1.2 0.128 ;
        RECT 1.198 0.346 1.2 0.3847 ;
        RECT 1.2 0.0427 1.232 0.0887 ;
        RECT 1.2 0.0887 1.232 0.1067 ;
        RECT 1.2 0.1067 1.232 0.128 ;
        RECT 1.2 0.346 1.232 0.3847 ;
        RECT 1.2 0.3847 1.232 0.3853 ;
        RECT 1.2 0.3853 1.232 0.4693 ;
        RECT 1.232 0.0887 1.266 0.1067 ;
        RECT 1.232 0.1067 1.266 0.128 ;
        RECT 1.232 0.346 1.266 0.3847 ;
        RECT 1.232 0.3847 1.266 0.3853 ;
        RECT 1.266 0.0887 1.294 0.1067 ;
        RECT 1.266 0.1067 1.294 0.128 ;
        RECT 1.266 0.128 1.294 0.346 ;
        RECT 1.266 0.346 1.294 0.3847 ;
        RECT 1.266 0.3847 1.294 0.3853 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.183 0.5307 ;
        RECT 1.183 0.4933 1.198 0.5307 ;
        RECT 1.198 0.4933 1.354 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.354 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2867 ;
        RECT 0.05 0.2867 0.078 0.4253 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.222 0.2267 ;
        RECT 0.178 0.2267 0.222 0.2867 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.37 0.0867 ;
        RECT 0.1533 0.1533 0.37 0.172 ;
        RECT 0.23 0.3827 0.37 0.4013 ;
        RECT 0.37 0.0679 0.398 0.0867 ;
        RECT 0.37 0.1533 0.398 0.172 ;
        RECT 0.37 0.172 0.398 0.1906 ;
        RECT 0.37 0.1906 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.3827 ;
        RECT 0.37 0.3827 0.398 0.4013 ;
        RECT 0.398 0.0679 0.6899 0.0867 ;
        RECT 0.6899 0.0679 0.718 0.0867 ;
        RECT 0.6899 0.0867 0.718 0.1533 ;
        RECT 0.6899 0.1533 0.718 0.172 ;
        RECT 0.6899 0.172 0.718 0.1906 ;
        RECT 0.6899 0.1906 0.718 0.228 ;
        RECT 0.718 0.172 1.198 0.1906 ;
        RECT 0.122 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.434 0.1293 ;
        RECT 0.274 0.4253 0.434 0.444 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.2573 ;
        RECT 0.434 0.2573 0.462 0.2687 ;
        RECT 0.434 0.2687 0.462 0.3073 ;
        RECT 0.434 0.3073 0.462 0.4253 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.4253 0.66 0.444 ;
        RECT 0.66 0.2573 0.718 0.2687 ;
        RECT 0.66 0.2687 0.718 0.3073 ;
        RECT 0.66 0.3073 0.718 0.4253 ;
        RECT 0.66 0.4253 0.718 0.444 ;
        RECT 0.718 0.2687 1.183 0.3073 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2867 ;
        RECT 0.05 0.2867 0.078 0.4253 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.222 0.2267 ;
        RECT 0.178 0.2267 0.222 0.2867 ;
        RECT 0.146 0.3827 0.202 0.4013 ;
        RECT 0.202 0.0679 0.23 0.0867 ;
        RECT 0.202 0.0867 0.1533 0.1533 ;
        RECT 0.202 0.1533 0.1533 0.172 ;
        RECT 0.202 0.3827 0.23 0.4013 ;
        RECT 0.23 0.0679 0.37 0.0867 ;
        RECT 0.1533 0.1533 0.37 0.172 ;
        RECT 0.23 0.3827 0.37 0.4013 ;
        RECT 0.37 0.0679 0.398 0.0867 ;
        RECT 0.37 0.1533 0.398 0.172 ;
        RECT 0.37 0.172 0.398 0.1906 ;
        RECT 0.37 0.1906 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.3827 ;
        RECT 0.37 0.3827 0.398 0.4013 ;
        RECT 0.398 0.0679 0.6899 0.0867 ;
        RECT 0.6899 0.0679 0.718 0.0867 ;
        RECT 0.6899 0.0867 0.718 0.1533 ;
        RECT 0.6899 0.1533 0.718 0.172 ;
        RECT 0.6899 0.172 0.718 0.1906 ;
        RECT 0.6899 0.1906 0.718 0.228 ;
        RECT 0.718 0.172 1.198 0.1906 ;
        RECT 0.122 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.434 0.1293 ;
        RECT 0.274 0.4253 0.434 0.444 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1293 0.462 0.2573 ;
        RECT 0.434 0.2573 0.462 0.2687 ;
        RECT 0.434 0.2687 0.462 0.3073 ;
        RECT 0.434 0.3073 0.462 0.4253 ;
        RECT 0.434 0.4253 0.462 0.444 ;
        RECT 0.462 0.4253 0.66 0.444 ;
        RECT 0.66 0.2573 0.718 0.2687 ;
        RECT 0.66 0.2687 0.718 0.3073 ;
        RECT 0.66 0.3073 0.718 0.4253 ;
        RECT 0.66 0.4253 0.718 0.444 ;
        RECT 0.718 0.2687 1.183 0.3073 ;
  END
END TBUF_X8_8T

MACRO TBUF_X12_8T
  CLASS core ;
  FOREIGN TBUF_X12_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.728 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.3587 ;
        RECT 0.1419 0.34 0.206 0.3587 ;
        RECT 0.206 0.34 0.242 0.3587 ;
        RECT 0.242 0.204 0.27 0.256 ;
        RECT 0.242 0.256 0.27 0.34 ;
        RECT 0.242 0.34 0.27 0.3587 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.268 0.498 0.2987 ;
        RECT 0.498 0.2306 0.526 0.268 ;
        RECT 0.498 0.268 0.526 0.2987 ;
        RECT 0.526 0.268 0.626 0.2987 ;
        RECT 0.626 0.268 0.654 0.2987 ;
        RECT 0.626 0.2987 0.654 0.384 ;
        RECT 0.654 0.268 0.71 0.2987 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.684 0.5307 ;
        RECT 1.684 0.4933 1.738 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 1.738 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2373 ;
        RECT 0.37 0.2373 0.398 0.252 ;
        RECT 0.37 0.252 0.398 0.284 ;
        RECT 0.37 0.284 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.783 0.444 ;
        RECT 0.783 0.2373 0.839 0.252 ;
        RECT 0.783 0.252 0.839 0.284 ;
        RECT 0.783 0.284 0.839 0.4253 ;
        RECT 0.783 0.4253 0.839 0.444 ;
        RECT 0.839 0.252 1.557 0.284 ;
        RECT 0.882 0.0679 0.931 0.0867 ;
        RECT 0.931 0.0679 0.989 0.0867 ;
        RECT 0.931 0.3547 0.989 0.3759 ;
        RECT 0.931 0.3759 0.989 0.4133 ;
        RECT 0.989 0.0679 1.572 0.0867 ;
        RECT 0.989 0.3547 1.572 0.3759 ;
        RECT 1.572 0.0487 1.586 0.0679 ;
        RECT 1.572 0.0679 1.586 0.0867 ;
        RECT 1.572 0.3547 1.586 0.3759 ;
        RECT 1.586 0.0487 1.614 0.0679 ;
        RECT 1.586 0.0679 1.614 0.0867 ;
        RECT 1.586 0.3547 1.614 0.3759 ;
        RECT 1.586 0.3759 1.614 0.4133 ;
        RECT 1.586 0.4133 1.614 0.41334 ;
        RECT 1.614 0.0487 1.6279 0.0679 ;
        RECT 1.614 0.0679 1.6279 0.0867 ;
        RECT 1.614 0.3547 1.6279 0.3759 ;
        RECT 1.6279 0.0679 1.629 0.0867 ;
        RECT 1.6279 0.3547 1.629 0.3759 ;
        RECT 1.629 0.0679 1.684 0.0867 ;
        RECT 1.629 0.0867 1.684 0.3547 ;
        RECT 1.629 0.3547 1.684 0.3759 ;
        RECT 0.05 0.1159 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.448 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.1419 0.0679 0.146 0.0867 ;
        RECT 0.1419 0.0867 0.146 0.1533 ;
        RECT 0.1419 0.1533 0.146 0.1667 ;
        RECT 0.1419 0.1667 0.146 0.16678 ;
        RECT 0.146 0.0679 0.17 0.0867 ;
        RECT 0.146 0.0867 0.17 0.1533 ;
        RECT 0.146 0.1533 0.17 0.1667 ;
        RECT 0.146 0.1667 0.17 0.16678 ;
        RECT 0.146 0.3827 0.17 0.4013 ;
        RECT 0.17 0.0679 0.306 0.0867 ;
        RECT 0.17 0.1533 0.306 0.1667 ;
        RECT 0.17 0.1667 0.306 0.16678 ;
        RECT 0.17 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.1667 ;
        RECT 0.306 0.1667 0.334 0.16678 ;
        RECT 0.306 0.172 0.334 0.196 ;
        RECT 0.306 0.196 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.782 0.0867 ;
        RECT 0.782 0.0679 0.8139 0.0867 ;
        RECT 0.782 0.0867 0.8139 0.1533 ;
        RECT 0.782 0.1533 0.8139 0.1667 ;
        RECT 0.782 0.1667 0.8139 0.16678 ;
        RECT 0.782 0.172 0.8139 0.196 ;
        RECT 0.8139 0.1667 1.593 0.16678 ;
        RECT 0.8139 0.172 1.593 0.196 ;
      LAYER M1 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.37 0.1293 ;
        RECT 0.274 0.4253 0.37 0.444 ;
        RECT 0.37 0.1107 0.398 0.1293 ;
        RECT 0.37 0.1293 0.398 0.2373 ;
        RECT 0.37 0.2373 0.398 0.252 ;
        RECT 0.37 0.252 0.398 0.284 ;
        RECT 0.37 0.284 0.398 0.4253 ;
        RECT 0.37 0.4253 0.398 0.444 ;
        RECT 0.398 0.4253 0.783 0.444 ;
        RECT 0.783 0.2373 0.839 0.252 ;
        RECT 0.783 0.252 0.839 0.284 ;
        RECT 0.783 0.284 0.839 0.4253 ;
        RECT 0.783 0.4253 0.839 0.444 ;
        RECT 0.839 0.252 1.557 0.284 ;
        RECT 0.882 0.0679 0.931 0.0867 ;
        RECT 0.931 0.0679 0.989 0.0867 ;
        RECT 0.931 0.3547 0.989 0.3759 ;
        RECT 0.931 0.3759 0.989 0.4133 ;
        RECT 0.989 0.0679 1.572 0.0867 ;
        RECT 0.989 0.3547 1.572 0.3759 ;
        RECT 1.572 0.0487 1.586 0.0679 ;
        RECT 1.572 0.0679 1.586 0.0867 ;
        RECT 1.572 0.3547 1.586 0.3759 ;
        RECT 1.586 0.0487 1.614 0.0679 ;
        RECT 1.586 0.0679 1.614 0.0867 ;
        RECT 1.586 0.3547 1.614 0.3759 ;
        RECT 1.586 0.3759 1.614 0.4133 ;
        RECT 1.586 0.4133 1.614 0.41334 ;
        RECT 1.614 0.0487 1.6279 0.0679 ;
        RECT 1.614 0.0679 1.6279 0.0867 ;
        RECT 1.614 0.3547 1.6279 0.3759 ;
        RECT 1.6279 0.0679 1.629 0.0867 ;
        RECT 1.6279 0.3547 1.629 0.3759 ;
        RECT 1.629 0.0679 1.684 0.0867 ;
        RECT 1.629 0.0867 1.684 0.3547 ;
        RECT 1.629 0.3547 1.684 0.3759 ;
        RECT 0.05 0.1159 0.078 0.208 ;
        RECT 0.05 0.208 0.078 0.2267 ;
        RECT 0.05 0.2267 0.078 0.2693 ;
        RECT 0.05 0.2693 0.078 0.448 ;
        RECT 0.078 0.208 0.178 0.2267 ;
        RECT 0.178 0.208 0.206 0.2267 ;
        RECT 0.178 0.2267 0.206 0.2693 ;
        RECT 0.1419 0.0679 0.146 0.0867 ;
        RECT 0.1419 0.0867 0.146 0.1533 ;
        RECT 0.1419 0.1533 0.146 0.1667 ;
        RECT 0.1419 0.1667 0.146 0.16678 ;
        RECT 0.146 0.0679 0.17 0.0867 ;
        RECT 0.146 0.0867 0.17 0.1533 ;
        RECT 0.146 0.1533 0.17 0.1667 ;
        RECT 0.146 0.1667 0.17 0.16678 ;
        RECT 0.146 0.3827 0.17 0.4013 ;
        RECT 0.17 0.0679 0.306 0.0867 ;
        RECT 0.17 0.1533 0.306 0.1667 ;
        RECT 0.17 0.1667 0.306 0.16678 ;
        RECT 0.17 0.3827 0.306 0.4013 ;
        RECT 0.306 0.0679 0.334 0.0867 ;
        RECT 0.306 0.1533 0.334 0.1667 ;
        RECT 0.306 0.1667 0.334 0.16678 ;
        RECT 0.306 0.172 0.334 0.196 ;
        RECT 0.306 0.196 0.334 0.3827 ;
        RECT 0.306 0.3827 0.334 0.4013 ;
        RECT 0.334 0.0679 0.782 0.0867 ;
        RECT 0.782 0.0679 0.8139 0.0867 ;
        RECT 0.782 0.0867 0.8139 0.1533 ;
        RECT 0.782 0.1533 0.8139 0.1667 ;
        RECT 0.782 0.1667 0.8139 0.16678 ;
        RECT 0.782 0.172 0.8139 0.196 ;
        RECT 0.8139 0.1667 1.593 0.16678 ;
        RECT 0.8139 0.172 1.593 0.196 ;
  END
END TBUF_X12_8T

MACRO TBUF_X16_8T
  CLASS core ;
  FOREIGN TBUF_X16_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.112 BY 0.512 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.26 0.1419 0.324 ;
        RECT 0.114 0.324 0.1419 0.3427 ;
        RECT 0.1419 0.324 0.1739 0.3427 ;
        RECT 0.1739 0.324 0.24 0.3427 ;
        RECT 0.24 0.2133 0.272 0.26 ;
        RECT 0.24 0.26 0.272 0.324 ;
        RECT 0.24 0.324 0.272 0.3427 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.462 0.268 0.562 0.2987 ;
        RECT 0.562 0.2306 0.59 0.268 ;
        RECT 0.562 0.268 0.59 0.2987 ;
        RECT 0.59 0.268 0.6899 0.2987 ;
        RECT 0.6899 0.268 0.718 0.2987 ;
        RECT 0.6899 0.2987 0.718 0.384 ;
        RECT 0.718 0.268 0.902 0.2987 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.0427 1.104 0.0946 ;
        RECT 1.072 0.0946 1.104 0.1333 ;
        RECT 1.072 0.3467 1.104 0.384 ;
        RECT 1.072 0.384 1.104 0.4693 ;
        RECT 1.104 0.0946 1.968 0.1333 ;
        RECT 1.104 0.3467 1.968 0.384 ;
        RECT 1.968 0.0427 1.98 0.0946 ;
        RECT 1.968 0.0946 1.98 0.1333 ;
        RECT 1.968 0.3467 1.98 0.384 ;
        RECT 1.968 0.384 1.98 0.4693 ;
        RECT 1.98 0.0427 1.998 0.0946 ;
        RECT 1.98 0.0946 1.998 0.1333 ;
        RECT 1.98 0.3467 1.998 0.384 ;
        RECT 1.98 0.384 1.998 0.4693 ;
        RECT 1.998 0.0427 2 0.0946 ;
        RECT 1.998 0.0946 2 0.1333 ;
        RECT 1.998 0.3467 2 0.384 ;
        RECT 1.998 0.384 2 0.4693 ;
        RECT 2 0.0946 2.0339 0.1333 ;
        RECT 2 0.3467 2.0339 0.384 ;
        RECT 2.0339 0.0946 2.062 0.1333 ;
        RECT 2.0339 0.1333 2.062 0.3467 ;
        RECT 2.0339 0.3467 2.062 0.384 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 1.98 0.5307 ;
        RECT 1.98 0.4933 1.998 0.5307 ;
        RECT 1.998 0.4933 2.122 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 2.122 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.1747 ;
        RECT 0.05 0.1747 0.078 0.1933 ;
        RECT 0.05 0.1933 0.078 0.2306 ;
        RECT 0.05 0.2306 0.078 0.4 ;
        RECT 0.078 0.1747 0.1419 0.1933 ;
        RECT 0.1419 0.1747 0.1739 0.1933 ;
        RECT 0.1419 0.1933 0.1739 0.2306 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.398 0.132 ;
        RECT 0.274 0.4253 0.398 0.444 ;
        RECT 0.398 0.1107 0.426 0.132 ;
        RECT 0.398 0.132 0.426 0.2687 ;
        RECT 0.398 0.2687 0.426 0.3073 ;
        RECT 0.398 0.3073 0.426 0.4253 ;
        RECT 0.398 0.4253 0.426 0.444 ;
        RECT 0.426 0.4253 0.946 0.444 ;
        RECT 0.946 0.2687 0.974 0.3073 ;
        RECT 0.946 0.3073 0.974 0.4253 ;
        RECT 0.946 0.4253 0.974 0.444 ;
        RECT 0.974 0.2687 1.98 0.3073 ;
        RECT 0.146 0.3786 0.21 0.4013 ;
        RECT 0.21 0.0679 0.238 0.0867 ;
        RECT 0.21 0.0867 0.238 0.156 ;
        RECT 0.21 0.156 0.238 0.1747 ;
        RECT 0.21 0.3786 0.238 0.4013 ;
        RECT 0.238 0.0679 0.326 0.0867 ;
        RECT 0.238 0.156 0.326 0.1747 ;
        RECT 0.238 0.3786 0.326 0.4013 ;
        RECT 0.326 0.0679 0.362 0.0867 ;
        RECT 0.326 0.156 0.362 0.1747 ;
        RECT 0.326 0.1747 0.362 0.182 ;
        RECT 0.326 0.182 0.362 0.2207 ;
        RECT 0.326 0.2207 0.362 0.3786 ;
        RECT 0.326 0.3786 0.362 0.4013 ;
        RECT 0.362 0.0679 0.946 0.0867 ;
        RECT 0.946 0.0679 0.974 0.0867 ;
        RECT 0.946 0.0867 0.974 0.156 ;
        RECT 0.946 0.156 0.974 0.1747 ;
        RECT 0.946 0.1747 0.974 0.182 ;
        RECT 0.946 0.182 0.974 0.2207 ;
        RECT 0.974 0.182 1.998 0.2207 ;
      LAYER M1 ;
        RECT 0.05 0.048 0.078 0.1747 ;
        RECT 0.05 0.1747 0.078 0.1933 ;
        RECT 0.05 0.1933 0.078 0.2306 ;
        RECT 0.05 0.2306 0.078 0.4 ;
        RECT 0.078 0.1747 0.1419 0.1933 ;
        RECT 0.1419 0.1747 0.1739 0.1933 ;
        RECT 0.1419 0.1933 0.1739 0.2306 ;
        RECT 0.146 0.4253 0.274 0.444 ;
        RECT 0.274 0.1107 0.398 0.132 ;
        RECT 0.274 0.4253 0.398 0.444 ;
        RECT 0.398 0.1107 0.426 0.132 ;
        RECT 0.398 0.132 0.426 0.2687 ;
        RECT 0.398 0.2687 0.426 0.3073 ;
        RECT 0.398 0.3073 0.426 0.4253 ;
        RECT 0.398 0.4253 0.426 0.444 ;
        RECT 0.426 0.4253 0.946 0.444 ;
        RECT 0.946 0.2687 0.974 0.3073 ;
        RECT 0.946 0.3073 0.974 0.4253 ;
        RECT 0.946 0.4253 0.974 0.444 ;
        RECT 0.974 0.2687 1.98 0.3073 ;
        RECT 0.146 0.3786 0.21 0.4013 ;
        RECT 0.21 0.0679 0.238 0.0867 ;
        RECT 0.21 0.0867 0.238 0.156 ;
        RECT 0.21 0.156 0.238 0.1747 ;
        RECT 0.21 0.3786 0.238 0.4013 ;
        RECT 0.238 0.0679 0.326 0.0867 ;
        RECT 0.238 0.156 0.326 0.1747 ;
        RECT 0.238 0.3786 0.326 0.4013 ;
        RECT 0.326 0.0679 0.362 0.0867 ;
        RECT 0.326 0.156 0.362 0.1747 ;
        RECT 0.326 0.1747 0.362 0.182 ;
        RECT 0.326 0.182 0.362 0.2207 ;
        RECT 0.326 0.2207 0.362 0.3786 ;
        RECT 0.326 0.3786 0.362 0.4013 ;
        RECT 0.362 0.0679 0.946 0.0867 ;
        RECT 0.946 0.0679 0.974 0.0867 ;
        RECT 0.946 0.0867 0.974 0.156 ;
        RECT 0.946 0.156 0.974 0.1747 ;
        RECT 0.946 0.1747 0.974 0.182 ;
        RECT 0.946 0.182 0.974 0.2207 ;
        RECT 0.974 0.182 1.998 0.2207 ;
  END
END TBUF_X16_8T

MACRO TIEH_8T
  CLASS core ;
  FOREIGN TIEH_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.3153 0.1419 0.4693 ;
        RECT 0.1419 0.3153 0.147 0.4693 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.286 ;
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.286 ;
  END
END TIEH_8T

MACRO TIEL_8T
  CLASS core ;
  FOREIGN TIEL_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.512 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.0427 0.147 0.1773 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.1419 0.5307 ;
        RECT 0.1419 0.4933 0.202 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.202 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.224 0.1419 0.448 ;
      LAYER M1 ;
        RECT 0.114 0.224 0.1419 0.448 ;
  END
END TIEL_8T

MACRO XNOR2_X1_8T
  CLASS core ;
  FOREIGN XNOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.168 0.21 0.1867 ;
        RECT 0.178 0.1867 0.21 0.2853 ;
        RECT 0.21 0.168 0.37 0.1867 ;
        RECT 0.37 0.168 0.398 0.1867 ;
        RECT 0.37 0.1867 0.398 0.2853 ;
        RECT 0.37 0.2853 0.398 0.2987 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.1613 0.078 0.2133 ;
        RECT 0.05 0.2133 0.078 0.4507 ;
        RECT 0.05 0.4507 0.078 0.4693 ;
        RECT 0.078 0.4507 0.274 0.4693 ;
        RECT 0.274 0.4507 0.498 0.4693 ;
        RECT 0.498 0.2133 0.526 0.4507 ;
        RECT 0.498 0.4507 0.526 0.4693 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.364 0.302 0.3647 ;
        RECT 0.278 0.3647 0.302 0.4007 ;
        RECT 0.278 0.4007 0.302 0.4013 ;
        RECT 0.302 0.1107 0.334 0.1293 ;
        RECT 0.302 0.364 0.334 0.3647 ;
        RECT 0.302 0.3647 0.334 0.4007 ;
        RECT 0.302 0.4007 0.334 0.4013 ;
        RECT 0.334 0.1107 0.434 0.1293 ;
        RECT 0.334 0.3647 0.434 0.4007 ;
        RECT 0.434 0.1107 0.462 0.1293 ;
        RECT 0.434 0.1653 0.462 0.184 ;
        RECT 0.434 0.184 0.462 0.364 ;
        RECT 0.434 0.364 0.462 0.3647 ;
        RECT 0.434 0.3647 0.462 0.4007 ;
        RECT 0.462 0.1107 0.493 0.1293 ;
        RECT 0.462 0.1653 0.493 0.184 ;
        RECT 0.493 0.1107 0.531 0.1293 ;
        RECT 0.493 0.1293 0.531 0.1653 ;
        RECT 0.493 0.1653 0.531 0.184 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.274 0.5307 ;
        RECT 0.274 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.0679 0.535 0.0867 ;
        RECT 0.114 0.1227 0.1419 0.144 ;
        RECT 0.114 0.144 0.1419 0.2267 ;
        RECT 0.114 0.2267 0.1419 0.3093 ;
        RECT 0.114 0.3093 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.368 ;
        RECT 0.1419 0.1227 0.234 0.144 ;
        RECT 0.1419 0.3093 0.234 0.328 ;
        RECT 0.234 0.3093 0.246 0.328 ;
        RECT 0.246 0.2267 0.274 0.3093 ;
        RECT 0.246 0.3093 0.274 0.328 ;
      LAYER M1 ;
        RECT 0.21 0.0679 0.535 0.0867 ;
        RECT 0.114 0.1227 0.1419 0.144 ;
        RECT 0.114 0.144 0.1419 0.2267 ;
        RECT 0.114 0.2267 0.1419 0.3093 ;
        RECT 0.114 0.3093 0.1419 0.328 ;
        RECT 0.114 0.328 0.1419 0.368 ;
        RECT 0.1419 0.1227 0.234 0.144 ;
        RECT 0.1419 0.3093 0.234 0.328 ;
        RECT 0.234 0.3093 0.246 0.328 ;
        RECT 0.246 0.2267 0.274 0.3093 ;
        RECT 0.246 0.3093 0.274 0.328 ;
  END
END XNOR2_X1_8T

MACRO XOR2_X1_8T
  CLASS core ;
  FOREIGN XOR2_X1_8T 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.512 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.2293 0.21 0.324 ;
        RECT 0.178 0.324 0.21 0.3427 ;
        RECT 0.21 0.324 0.274 0.3427 ;
        RECT 0.274 0.324 0.37 0.3427 ;
        RECT 0.37 0.2133 0.398 0.2293 ;
        RECT 0.37 0.2293 0.398 0.324 ;
        RECT 0.37 0.324 0.398 0.3427 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.0427 0.078 0.0613 ;
        RECT 0.05 0.0613 0.078 0.2987 ;
        RECT 0.05 0.2987 0.078 0.3507 ;
        RECT 0.078 0.0427 0.498 0.0613 ;
        RECT 0.498 0.0427 0.526 0.0613 ;
        RECT 0.498 0.0613 0.526 0.2987 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.275 0.1087 0.315 0.1093 ;
        RECT 0.275 0.1093 0.315 0.148 ;
        RECT 0.315 0.1087 0.334 0.1093 ;
        RECT 0.315 0.1093 0.334 0.148 ;
        RECT 0.315 0.3827 0.334 0.4013 ;
        RECT 0.334 0.1093 0.434 0.148 ;
        RECT 0.334 0.3827 0.434 0.4013 ;
        RECT 0.434 0.1093 0.462 0.148 ;
        RECT 0.434 0.148 0.462 0.328 ;
        RECT 0.434 0.328 0.462 0.3467 ;
        RECT 0.434 0.3827 0.462 0.4013 ;
        RECT 0.462 0.328 0.496 0.3467 ;
        RECT 0.462 0.3827 0.496 0.4013 ;
        RECT 0.496 0.328 0.34678 0.3467 ;
        RECT 0.496 0.3467 0.34678 0.3827 ;
        RECT 0.496 0.3827 0.528 0.4013 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.4933 0.535 0.5307 ;
        RECT 0.535 0.4933 0.586 0.5307 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.0187 0.586 0.0187 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.246 0.4253 0.535 0.444 ;
        RECT 0.114 0.0907 0.1419 0.1867 ;
        RECT 0.114 0.1867 0.1419 0.2053 ;
        RECT 0.114 0.2053 0.1419 0.288 ;
        RECT 0.114 0.288 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.3893 ;
        RECT 0.1419 0.1867 0.246 0.2053 ;
        RECT 0.1419 0.368 0.246 0.3893 ;
        RECT 0.246 0.1867 0.247 0.2053 ;
        RECT 0.246 0.2053 0.247 0.288 ;
        RECT 0.246 0.368 0.247 0.3893 ;
        RECT 0.247 0.1867 0.274 0.2053 ;
        RECT 0.247 0.2053 0.274 0.288 ;
      LAYER M1 ;
        RECT 0.246 0.4253 0.535 0.444 ;
        RECT 0.114 0.0907 0.1419 0.1867 ;
        RECT 0.114 0.1867 0.1419 0.2053 ;
        RECT 0.114 0.2053 0.1419 0.288 ;
        RECT 0.114 0.288 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.3893 ;
        RECT 0.1419 0.1867 0.246 0.2053 ;
        RECT 0.1419 0.368 0.246 0.3893 ;
        RECT 0.246 0.1867 0.247 0.2053 ;
        RECT 0.246 0.2053 0.247 0.288 ;
        RECT 0.246 0.368 0.247 0.3893 ;
        RECT 0.247 0.1867 0.274 0.2053 ;
        RECT 0.247 0.2053 0.274 0.288 ;
  END
END XOR2_X1_8T

END LIBRARY
#
# End of file
#
